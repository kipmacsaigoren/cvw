///////////////////////////////////////////
// clmul.sv
//
// Written: Kevin Kim <kekim@hmc.edu> and Kip Macsai-Goren <kmacsaigoren@hmc.edu>
// Created: 1 February 2023
// Modified: 
//
// Purpose: Carry-Less multiplication unit
//
// Documentation: RISC-V System on Chip Design Chapter 15
// 
// A component of the CORE-V-WALLY configurable RISC-V project.
// 
// Copyright (C) 2021-23 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`include "wally-config.vh"

module clmulopt #(parameter WIDTH=32) (
  input  logic [WIDTH-1:0] X, Y,             // Operands
  output logic [WIDTH-1:0] ClmulResult);     // ZBS result

  if (WIDTH == 64) begin
    assign S0 = X[0] & Y[0];
    assign ClmulResult[0] = S0;
    assign S64 = X[0] & Y[1];
    assign S65 = (X[1] & Y[0]) ^ S64;
    assign ClmulResult[1] = S65;
    assign S128 = X[0] & Y[2];
    assign S129 = (X[1] & Y[1]) ^ S128;
    assign S130 = (X[2] & Y[0]) ^ S129;
    assign ClmulResult[2] = S130;
    assign S192 = X[0] & Y[3];
    assign S193 = (X[1] & Y[2]) ^ S192;
    assign S194 = (X[2] & Y[1]) ^ S193;
    assign S195 = (X[3] & Y[0]) ^ S194;
    assign ClmulResult[3] = S195;
    assign S256 = X[0] & Y[4];
    assign S257 = (X[1] & Y[3]) ^ S256;
    assign S258 = (X[2] & Y[2]) ^ S257;
    assign S259 = (X[3] & Y[1]) ^ S258;
    assign S260 = (X[4] & Y[0]) ^ S259;
    assign ClmulResult[4] = S260;
    assign S320 = X[0] & Y[5];
    assign S321 = (X[1] & Y[4]) ^ S320;
    assign S322 = (X[2] & Y[3]) ^ S321;
    assign S323 = (X[3] & Y[2]) ^ S322;
    assign S324 = (X[4] & Y[1]) ^ S323;
    assign S325 = (X[5] & Y[0]) ^ S324;
    assign ClmulResult[5] = S325;
    assign S384 = X[0] & Y[6];
    assign S385 = (X[1] & Y[5]) ^ S384;
    assign S386 = (X[2] & Y[4]) ^ S385;
    assign S387 = (X[3] & Y[3]) ^ S386;
    assign S388 = (X[4] & Y[2]) ^ S387;
    assign S389 = (X[5] & Y[1]) ^ S388;
    assign S390 = (X[6] & Y[0]) ^ S389;
    assign ClmulResult[6] = S390;
    assign S448 = X[0] & Y[7];
    assign S449 = (X[1] & Y[6]) ^ S448;
    assign S450 = (X[2] & Y[5]) ^ S449;
    assign S451 = (X[3] & Y[4]) ^ S450;
    assign S452 = (X[4] & Y[3]) ^ S451;
    assign S453 = (X[5] & Y[2]) ^ S452;
    assign S454 = (X[6] & Y[1]) ^ S453;
    assign S455 = (X[7] & Y[0]) ^ S454;
    assign ClmulResult[7] = S455;
    assign S512 = X[0] & Y[8];
    assign S513 = (X[1] & Y[7]) ^ S512;
    assign S514 = (X[2] & Y[6]) ^ S513;
    assign S515 = (X[3] & Y[5]) ^ S514;
    assign S516 = (X[4] & Y[4]) ^ S515;
    assign S517 = (X[5] & Y[3]) ^ S516;
    assign S518 = (X[6] & Y[2]) ^ S517;
    assign S519 = (X[7] & Y[1]) ^ S518;
    assign S520 = (X[8] & Y[0]) ^ S519;
    assign ClmulResult[8] = S520;
    assign S576 = X[0] & Y[9];
    assign S577 = (X[1] & Y[8]) ^ S576;
    assign S578 = (X[2] & Y[7]) ^ S577;
    assign S579 = (X[3] & Y[6]) ^ S578;
    assign S580 = (X[4] & Y[5]) ^ S579;
    assign S581 = (X[5] & Y[4]) ^ S580;
    assign S582 = (X[6] & Y[3]) ^ S581;
    assign S583 = (X[7] & Y[2]) ^ S582;
    assign S584 = (X[8] & Y[1]) ^ S583;
    assign S585 = (X[9] & Y[0]) ^ S584;
    assign ClmulResult[9] = S585;
    assign S640 = X[0] & Y[10];
    assign S641 = (X[1] & Y[9]) ^ S640;
    assign S642 = (X[2] & Y[8]) ^ S641;
    assign S643 = (X[3] & Y[7]) ^ S642;
    assign S644 = (X[4] & Y[6]) ^ S643;
    assign S645 = (X[5] & Y[5]) ^ S644;
    assign S646 = (X[6] & Y[4]) ^ S645;
    assign S647 = (X[7] & Y[3]) ^ S646;
    assign S648 = (X[8] & Y[2]) ^ S647;
    assign S649 = (X[9] & Y[1]) ^ S648;
    assign S650 = (X[10] & Y[0]) ^ S649;
    assign ClmulResult[10] = S650;
    assign S704 = X[0] & Y[11];
    assign S705 = (X[1] & Y[10]) ^ S704;
    assign S706 = (X[2] & Y[9]) ^ S705;
    assign S707 = (X[3] & Y[8]) ^ S706;
    assign S708 = (X[4] & Y[7]) ^ S707;
    assign S709 = (X[5] & Y[6]) ^ S708;
    assign S710 = (X[6] & Y[5]) ^ S709;
    assign S711 = (X[7] & Y[4]) ^ S710;
    assign S712 = (X[8] & Y[3]) ^ S711;
    assign S713 = (X[9] & Y[2]) ^ S712;
    assign S714 = (X[10] & Y[1]) ^ S713;
    assign S715 = (X[11] & Y[0]) ^ S714;
    assign ClmulResult[11] = S715;
    assign S768 = X[0] & Y[12];
    assign S769 = (X[1] & Y[11]) ^ S768;
    assign S770 = (X[2] & Y[10]) ^ S769;
    assign S771 = (X[3] & Y[9]) ^ S770;
    assign S772 = (X[4] & Y[8]) ^ S771;
    assign S773 = (X[5] & Y[7]) ^ S772;
    assign S774 = (X[6] & Y[6]) ^ S773;
    assign S775 = (X[7] & Y[5]) ^ S774;
    assign S776 = (X[8] & Y[4]) ^ S775;
    assign S777 = (X[9] & Y[3]) ^ S776;
    assign S778 = (X[10] & Y[2]) ^ S777;
    assign S779 = (X[11] & Y[1]) ^ S778;
    assign S780 = (X[12] & Y[0]) ^ S779;
    assign ClmulResult[12] = S780;
    assign S832 = X[0] & Y[13];
    assign S833 = (X[1] & Y[12]) ^ S832;
    assign S834 = (X[2] & Y[11]) ^ S833;
    assign S835 = (X[3] & Y[10]) ^ S834;
    assign S836 = (X[4] & Y[9]) ^ S835;
    assign S837 = (X[5] & Y[8]) ^ S836;
    assign S838 = (X[6] & Y[7]) ^ S837;
    assign S839 = (X[7] & Y[6]) ^ S838;
    assign S840 = (X[8] & Y[5]) ^ S839;
    assign S841 = (X[9] & Y[4]) ^ S840;
    assign S842 = (X[10] & Y[3]) ^ S841;
    assign S843 = (X[11] & Y[2]) ^ S842;
    assign S844 = (X[12] & Y[1]) ^ S843;
    assign S845 = (X[13] & Y[0]) ^ S844;
    assign ClmulResult[13] = S845;
    assign S896 = X[0] & Y[14];
    assign S897 = (X[1] & Y[13]) ^ S896;
    assign S898 = (X[2] & Y[12]) ^ S897;
    assign S899 = (X[3] & Y[11]) ^ S898;
    assign S900 = (X[4] & Y[10]) ^ S899;
    assign S901 = (X[5] & Y[9]) ^ S900;
    assign S902 = (X[6] & Y[8]) ^ S901;
    assign S903 = (X[7] & Y[7]) ^ S902;
    assign S904 = (X[8] & Y[6]) ^ S903;
    assign S905 = (X[9] & Y[5]) ^ S904;
    assign S906 = (X[10] & Y[4]) ^ S905;
    assign S907 = (X[11] & Y[3]) ^ S906;
    assign S908 = (X[12] & Y[2]) ^ S907;
    assign S909 = (X[13] & Y[1]) ^ S908;
    assign S910 = (X[14] & Y[0]) ^ S909;
    assign ClmulResult[14] = S910;
    assign S960 = X[0] & Y[15];
    assign S961 = (X[1] & Y[14]) ^ S960;
    assign S962 = (X[2] & Y[13]) ^ S961;
    assign S963 = (X[3] & Y[12]) ^ S962;
    assign S964 = (X[4] & Y[11]) ^ S963;
    assign S965 = (X[5] & Y[10]) ^ S964;
    assign S966 = (X[6] & Y[9]) ^ S965;
    assign S967 = (X[7] & Y[8]) ^ S966;
    assign S968 = (X[8] & Y[7]) ^ S967;
    assign S969 = (X[9] & Y[6]) ^ S968;
    assign S970 = (X[10] & Y[5]) ^ S969;
    assign S971 = (X[11] & Y[4]) ^ S970;
    assign S972 = (X[12] & Y[3]) ^ S971;
    assign S973 = (X[13] & Y[2]) ^ S972;
    assign S974 = (X[14] & Y[1]) ^ S973;
    assign S975 = (X[15] & Y[0]) ^ S974;
    assign ClmulResult[15] = S975;
    assign S1024 = X[0] & Y[16];
    assign S1025 = (X[1] & Y[15]) ^ S1024;
    assign S1026 = (X[2] & Y[14]) ^ S1025;
    assign S1027 = (X[3] & Y[13]) ^ S1026;
    assign S1028 = (X[4] & Y[12]) ^ S1027;
    assign S1029 = (X[5] & Y[11]) ^ S1028;
    assign S1030 = (X[6] & Y[10]) ^ S1029;
    assign S1031 = (X[7] & Y[9]) ^ S1030;
    assign S1032 = (X[8] & Y[8]) ^ S1031;
    assign S1033 = (X[9] & Y[7]) ^ S1032;
    assign S1034 = (X[10] & Y[6]) ^ S1033;
    assign S1035 = (X[11] & Y[5]) ^ S1034;
    assign S1036 = (X[12] & Y[4]) ^ S1035;
    assign S1037 = (X[13] & Y[3]) ^ S1036;
    assign S1038 = (X[14] & Y[2]) ^ S1037;
    assign S1039 = (X[15] & Y[1]) ^ S1038;
    assign S1040 = (X[16] & Y[0]) ^ S1039;
    assign ClmulResult[16] = S1040;
    assign S1088 = X[0] & Y[17];
    assign S1089 = (X[1] & Y[16]) ^ S1088;
    assign S1090 = (X[2] & Y[15]) ^ S1089;
    assign S1091 = (X[3] & Y[14]) ^ S1090;
    assign S1092 = (X[4] & Y[13]) ^ S1091;
    assign S1093 = (X[5] & Y[12]) ^ S1092;
    assign S1094 = (X[6] & Y[11]) ^ S1093;
    assign S1095 = (X[7] & Y[10]) ^ S1094;
    assign S1096 = (X[8] & Y[9]) ^ S1095;
    assign S1097 = (X[9] & Y[8]) ^ S1096;
    assign S1098 = (X[10] & Y[7]) ^ S1097;
    assign S1099 = (X[11] & Y[6]) ^ S1098;
    assign S1100 = (X[12] & Y[5]) ^ S1099;
    assign S1101 = (X[13] & Y[4]) ^ S1100;
    assign S1102 = (X[14] & Y[3]) ^ S1101;
    assign S1103 = (X[15] & Y[2]) ^ S1102;
    assign S1104 = (X[16] & Y[1]) ^ S1103;
    assign S1105 = (X[17] & Y[0]) ^ S1104;
    assign ClmulResult[17] = S1105;
    assign S1152 = X[0] & Y[18];
    assign S1153 = (X[1] & Y[17]) ^ S1152;
    assign S1154 = (X[2] & Y[16]) ^ S1153;
    assign S1155 = (X[3] & Y[15]) ^ S1154;
    assign S1156 = (X[4] & Y[14]) ^ S1155;
    assign S1157 = (X[5] & Y[13]) ^ S1156;
    assign S1158 = (X[6] & Y[12]) ^ S1157;
    assign S1159 = (X[7] & Y[11]) ^ S1158;
    assign S1160 = (X[8] & Y[10]) ^ S1159;
    assign S1161 = (X[9] & Y[9]) ^ S1160;
    assign S1162 = (X[10] & Y[8]) ^ S1161;
    assign S1163 = (X[11] & Y[7]) ^ S1162;
    assign S1164 = (X[12] & Y[6]) ^ S1163;
    assign S1165 = (X[13] & Y[5]) ^ S1164;
    assign S1166 = (X[14] & Y[4]) ^ S1165;
    assign S1167 = (X[15] & Y[3]) ^ S1166;
    assign S1168 = (X[16] & Y[2]) ^ S1167;
    assign S1169 = (X[17] & Y[1]) ^ S1168;
    assign S1170 = (X[18] & Y[0]) ^ S1169;
    assign ClmulResult[18] = S1170;
    assign S1216 = X[0] & Y[19];
    assign S1217 = (X[1] & Y[18]) ^ S1216;
    assign S1218 = (X[2] & Y[17]) ^ S1217;
    assign S1219 = (X[3] & Y[16]) ^ S1218;
    assign S1220 = (X[4] & Y[15]) ^ S1219;
    assign S1221 = (X[5] & Y[14]) ^ S1220;
    assign S1222 = (X[6] & Y[13]) ^ S1221;
    assign S1223 = (X[7] & Y[12]) ^ S1222;
    assign S1224 = (X[8] & Y[11]) ^ S1223;
    assign S1225 = (X[9] & Y[10]) ^ S1224;
    assign S1226 = (X[10] & Y[9]) ^ S1225;
    assign S1227 = (X[11] & Y[8]) ^ S1226;
    assign S1228 = (X[12] & Y[7]) ^ S1227;
    assign S1229 = (X[13] & Y[6]) ^ S1228;
    assign S1230 = (X[14] & Y[5]) ^ S1229;
    assign S1231 = (X[15] & Y[4]) ^ S1230;
    assign S1232 = (X[16] & Y[3]) ^ S1231;
    assign S1233 = (X[17] & Y[2]) ^ S1232;
    assign S1234 = (X[18] & Y[1]) ^ S1233;
    assign S1235 = (X[19] & Y[0]) ^ S1234;
    assign ClmulResult[19] = S1235;
    assign S1280 = X[0] & Y[20];
    assign S1281 = (X[1] & Y[19]) ^ S1280;
    assign S1282 = (X[2] & Y[18]) ^ S1281;
    assign S1283 = (X[3] & Y[17]) ^ S1282;
    assign S1284 = (X[4] & Y[16]) ^ S1283;
    assign S1285 = (X[5] & Y[15]) ^ S1284;
    assign S1286 = (X[6] & Y[14]) ^ S1285;
    assign S1287 = (X[7] & Y[13]) ^ S1286;
    assign S1288 = (X[8] & Y[12]) ^ S1287;
    assign S1289 = (X[9] & Y[11]) ^ S1288;
    assign S1290 = (X[10] & Y[10]) ^ S1289;
    assign S1291 = (X[11] & Y[9]) ^ S1290;
    assign S1292 = (X[12] & Y[8]) ^ S1291;
    assign S1293 = (X[13] & Y[7]) ^ S1292;
    assign S1294 = (X[14] & Y[6]) ^ S1293;
    assign S1295 = (X[15] & Y[5]) ^ S1294;
    assign S1296 = (X[16] & Y[4]) ^ S1295;
    assign S1297 = (X[17] & Y[3]) ^ S1296;
    assign S1298 = (X[18] & Y[2]) ^ S1297;
    assign S1299 = (X[19] & Y[1]) ^ S1298;
    assign S1300 = (X[20] & Y[0]) ^ S1299;
    assign ClmulResult[20] = S1300;
    assign S1344 = X[0] & Y[21];
    assign S1345 = (X[1] & Y[20]) ^ S1344;
    assign S1346 = (X[2] & Y[19]) ^ S1345;
    assign S1347 = (X[3] & Y[18]) ^ S1346;
    assign S1348 = (X[4] & Y[17]) ^ S1347;
    assign S1349 = (X[5] & Y[16]) ^ S1348;
    assign S1350 = (X[6] & Y[15]) ^ S1349;
    assign S1351 = (X[7] & Y[14]) ^ S1350;
    assign S1352 = (X[8] & Y[13]) ^ S1351;
    assign S1353 = (X[9] & Y[12]) ^ S1352;
    assign S1354 = (X[10] & Y[11]) ^ S1353;
    assign S1355 = (X[11] & Y[10]) ^ S1354;
    assign S1356 = (X[12] & Y[9]) ^ S1355;
    assign S1357 = (X[13] & Y[8]) ^ S1356;
    assign S1358 = (X[14] & Y[7]) ^ S1357;
    assign S1359 = (X[15] & Y[6]) ^ S1358;
    assign S1360 = (X[16] & Y[5]) ^ S1359;
    assign S1361 = (X[17] & Y[4]) ^ S1360;
    assign S1362 = (X[18] & Y[3]) ^ S1361;
    assign S1363 = (X[19] & Y[2]) ^ S1362;
    assign S1364 = (X[20] & Y[1]) ^ S1363;
    assign S1365 = (X[21] & Y[0]) ^ S1364;
    assign ClmulResult[21] = S1365;
    assign S1408 = X[0] & Y[22];
    assign S1409 = (X[1] & Y[21]) ^ S1408;
    assign S1410 = (X[2] & Y[20]) ^ S1409;
    assign S1411 = (X[3] & Y[19]) ^ S1410;
    assign S1412 = (X[4] & Y[18]) ^ S1411;
    assign S1413 = (X[5] & Y[17]) ^ S1412;
    assign S1414 = (X[6] & Y[16]) ^ S1413;
    assign S1415 = (X[7] & Y[15]) ^ S1414;
    assign S1416 = (X[8] & Y[14]) ^ S1415;
    assign S1417 = (X[9] & Y[13]) ^ S1416;
    assign S1418 = (X[10] & Y[12]) ^ S1417;
    assign S1419 = (X[11] & Y[11]) ^ S1418;
    assign S1420 = (X[12] & Y[10]) ^ S1419;
    assign S1421 = (X[13] & Y[9]) ^ S1420;
    assign S1422 = (X[14] & Y[8]) ^ S1421;
    assign S1423 = (X[15] & Y[7]) ^ S1422;
    assign S1424 = (X[16] & Y[6]) ^ S1423;
    assign S1425 = (X[17] & Y[5]) ^ S1424;
    assign S1426 = (X[18] & Y[4]) ^ S1425;
    assign S1427 = (X[19] & Y[3]) ^ S1426;
    assign S1428 = (X[20] & Y[2]) ^ S1427;
    assign S1429 = (X[21] & Y[1]) ^ S1428;
    assign S1430 = (X[22] & Y[0]) ^ S1429;
    assign ClmulResult[22] = S1430;
    assign S1472 = X[0] & Y[23];
    assign S1473 = (X[1] & Y[22]) ^ S1472;
    assign S1474 = (X[2] & Y[21]) ^ S1473;
    assign S1475 = (X[3] & Y[20]) ^ S1474;
    assign S1476 = (X[4] & Y[19]) ^ S1475;
    assign S1477 = (X[5] & Y[18]) ^ S1476;
    assign S1478 = (X[6] & Y[17]) ^ S1477;
    assign S1479 = (X[7] & Y[16]) ^ S1478;
    assign S1480 = (X[8] & Y[15]) ^ S1479;
    assign S1481 = (X[9] & Y[14]) ^ S1480;
    assign S1482 = (X[10] & Y[13]) ^ S1481;
    assign S1483 = (X[11] & Y[12]) ^ S1482;
    assign S1484 = (X[12] & Y[11]) ^ S1483;
    assign S1485 = (X[13] & Y[10]) ^ S1484;
    assign S1486 = (X[14] & Y[9]) ^ S1485;
    assign S1487 = (X[15] & Y[8]) ^ S1486;
    assign S1488 = (X[16] & Y[7]) ^ S1487;
    assign S1489 = (X[17] & Y[6]) ^ S1488;
    assign S1490 = (X[18] & Y[5]) ^ S1489;
    assign S1491 = (X[19] & Y[4]) ^ S1490;
    assign S1492 = (X[20] & Y[3]) ^ S1491;
    assign S1493 = (X[21] & Y[2]) ^ S1492;
    assign S1494 = (X[22] & Y[1]) ^ S1493;
    assign S1495 = (X[23] & Y[0]) ^ S1494;
    assign ClmulResult[23] = S1495;
    assign S1536 = X[0] & Y[24];
    assign S1537 = (X[1] & Y[23]) ^ S1536;
    assign S1538 = (X[2] & Y[22]) ^ S1537;
    assign S1539 = (X[3] & Y[21]) ^ S1538;
    assign S1540 = (X[4] & Y[20]) ^ S1539;
    assign S1541 = (X[5] & Y[19]) ^ S1540;
    assign S1542 = (X[6] & Y[18]) ^ S1541;
    assign S1543 = (X[7] & Y[17]) ^ S1542;
    assign S1544 = (X[8] & Y[16]) ^ S1543;
    assign S1545 = (X[9] & Y[15]) ^ S1544;
    assign S1546 = (X[10] & Y[14]) ^ S1545;
    assign S1547 = (X[11] & Y[13]) ^ S1546;
    assign S1548 = (X[12] & Y[12]) ^ S1547;
    assign S1549 = (X[13] & Y[11]) ^ S1548;
    assign S1550 = (X[14] & Y[10]) ^ S1549;
    assign S1551 = (X[15] & Y[9]) ^ S1550;
    assign S1552 = (X[16] & Y[8]) ^ S1551;
    assign S1553 = (X[17] & Y[7]) ^ S1552;
    assign S1554 = (X[18] & Y[6]) ^ S1553;
    assign S1555 = (X[19] & Y[5]) ^ S1554;
    assign S1556 = (X[20] & Y[4]) ^ S1555;
    assign S1557 = (X[21] & Y[3]) ^ S1556;
    assign S1558 = (X[22] & Y[2]) ^ S1557;
    assign S1559 = (X[23] & Y[1]) ^ S1558;
    assign S1560 = (X[24] & Y[0]) ^ S1559;
    assign ClmulResult[24] = S1560;
    assign S1600 = X[0] & Y[25];
    assign S1601 = (X[1] & Y[24]) ^ S1600;
    assign S1602 = (X[2] & Y[23]) ^ S1601;
    assign S1603 = (X[3] & Y[22]) ^ S1602;
    assign S1604 = (X[4] & Y[21]) ^ S1603;
    assign S1605 = (X[5] & Y[20]) ^ S1604;
    assign S1606 = (X[6] & Y[19]) ^ S1605;
    assign S1607 = (X[7] & Y[18]) ^ S1606;
    assign S1608 = (X[8] & Y[17]) ^ S1607;
    assign S1609 = (X[9] & Y[16]) ^ S1608;
    assign S1610 = (X[10] & Y[15]) ^ S1609;
    assign S1611 = (X[11] & Y[14]) ^ S1610;
    assign S1612 = (X[12] & Y[13]) ^ S1611;
    assign S1613 = (X[13] & Y[12]) ^ S1612;
    assign S1614 = (X[14] & Y[11]) ^ S1613;
    assign S1615 = (X[15] & Y[10]) ^ S1614;
    assign S1616 = (X[16] & Y[9]) ^ S1615;
    assign S1617 = (X[17] & Y[8]) ^ S1616;
    assign S1618 = (X[18] & Y[7]) ^ S1617;
    assign S1619 = (X[19] & Y[6]) ^ S1618;
    assign S1620 = (X[20] & Y[5]) ^ S1619;
    assign S1621 = (X[21] & Y[4]) ^ S1620;
    assign S1622 = (X[22] & Y[3]) ^ S1621;
    assign S1623 = (X[23] & Y[2]) ^ S1622;
    assign S1624 = (X[24] & Y[1]) ^ S1623;
    assign S1625 = (X[25] & Y[0]) ^ S1624;
    assign ClmulResult[25] = S1625;
    assign S1664 = X[0] & Y[26];
    assign S1665 = (X[1] & Y[25]) ^ S1664;
    assign S1666 = (X[2] & Y[24]) ^ S1665;
    assign S1667 = (X[3] & Y[23]) ^ S1666;
    assign S1668 = (X[4] & Y[22]) ^ S1667;
    assign S1669 = (X[5] & Y[21]) ^ S1668;
    assign S1670 = (X[6] & Y[20]) ^ S1669;
    assign S1671 = (X[7] & Y[19]) ^ S1670;
    assign S1672 = (X[8] & Y[18]) ^ S1671;
    assign S1673 = (X[9] & Y[17]) ^ S1672;
    assign S1674 = (X[10] & Y[16]) ^ S1673;
    assign S1675 = (X[11] & Y[15]) ^ S1674;
    assign S1676 = (X[12] & Y[14]) ^ S1675;
    assign S1677 = (X[13] & Y[13]) ^ S1676;
    assign S1678 = (X[14] & Y[12]) ^ S1677;
    assign S1679 = (X[15] & Y[11]) ^ S1678;
    assign S1680 = (X[16] & Y[10]) ^ S1679;
    assign S1681 = (X[17] & Y[9]) ^ S1680;
    assign S1682 = (X[18] & Y[8]) ^ S1681;
    assign S1683 = (X[19] & Y[7]) ^ S1682;
    assign S1684 = (X[20] & Y[6]) ^ S1683;
    assign S1685 = (X[21] & Y[5]) ^ S1684;
    assign S1686 = (X[22] & Y[4]) ^ S1685;
    assign S1687 = (X[23] & Y[3]) ^ S1686;
    assign S1688 = (X[24] & Y[2]) ^ S1687;
    assign S1689 = (X[25] & Y[1]) ^ S1688;
    assign S1690 = (X[26] & Y[0]) ^ S1689;
    assign ClmulResult[26] = S1690;
    assign S1728 = X[0] & Y[27];
    assign S1729 = (X[1] & Y[26]) ^ S1728;
    assign S1730 = (X[2] & Y[25]) ^ S1729;
    assign S1731 = (X[3] & Y[24]) ^ S1730;
    assign S1732 = (X[4] & Y[23]) ^ S1731;
    assign S1733 = (X[5] & Y[22]) ^ S1732;
    assign S1734 = (X[6] & Y[21]) ^ S1733;
    assign S1735 = (X[7] & Y[20]) ^ S1734;
    assign S1736 = (X[8] & Y[19]) ^ S1735;
    assign S1737 = (X[9] & Y[18]) ^ S1736;
    assign S1738 = (X[10] & Y[17]) ^ S1737;
    assign S1739 = (X[11] & Y[16]) ^ S1738;
    assign S1740 = (X[12] & Y[15]) ^ S1739;
    assign S1741 = (X[13] & Y[14]) ^ S1740;
    assign S1742 = (X[14] & Y[13]) ^ S1741;
    assign S1743 = (X[15] & Y[12]) ^ S1742;
    assign S1744 = (X[16] & Y[11]) ^ S1743;
    assign S1745 = (X[17] & Y[10]) ^ S1744;
    assign S1746 = (X[18] & Y[9]) ^ S1745;
    assign S1747 = (X[19] & Y[8]) ^ S1746;
    assign S1748 = (X[20] & Y[7]) ^ S1747;
    assign S1749 = (X[21] & Y[6]) ^ S1748;
    assign S1750 = (X[22] & Y[5]) ^ S1749;
    assign S1751 = (X[23] & Y[4]) ^ S1750;
    assign S1752 = (X[24] & Y[3]) ^ S1751;
    assign S1753 = (X[25] & Y[2]) ^ S1752;
    assign S1754 = (X[26] & Y[1]) ^ S1753;
    assign S1755 = (X[27] & Y[0]) ^ S1754;
    assign ClmulResult[27] = S1755;
    assign S1792 = X[0] & Y[28];
    assign S1793 = (X[1] & Y[27]) ^ S1792;
    assign S1794 = (X[2] & Y[26]) ^ S1793;
    assign S1795 = (X[3] & Y[25]) ^ S1794;
    assign S1796 = (X[4] & Y[24]) ^ S1795;
    assign S1797 = (X[5] & Y[23]) ^ S1796;
    assign S1798 = (X[6] & Y[22]) ^ S1797;
    assign S1799 = (X[7] & Y[21]) ^ S1798;
    assign S1800 = (X[8] & Y[20]) ^ S1799;
    assign S1801 = (X[9] & Y[19]) ^ S1800;
    assign S1802 = (X[10] & Y[18]) ^ S1801;
    assign S1803 = (X[11] & Y[17]) ^ S1802;
    assign S1804 = (X[12] & Y[16]) ^ S1803;
    assign S1805 = (X[13] & Y[15]) ^ S1804;
    assign S1806 = (X[14] & Y[14]) ^ S1805;
    assign S1807 = (X[15] & Y[13]) ^ S1806;
    assign S1808 = (X[16] & Y[12]) ^ S1807;
    assign S1809 = (X[17] & Y[11]) ^ S1808;
    assign S1810 = (X[18] & Y[10]) ^ S1809;
    assign S1811 = (X[19] & Y[9]) ^ S1810;
    assign S1812 = (X[20] & Y[8]) ^ S1811;
    assign S1813 = (X[21] & Y[7]) ^ S1812;
    assign S1814 = (X[22] & Y[6]) ^ S1813;
    assign S1815 = (X[23] & Y[5]) ^ S1814;
    assign S1816 = (X[24] & Y[4]) ^ S1815;
    assign S1817 = (X[25] & Y[3]) ^ S1816;
    assign S1818 = (X[26] & Y[2]) ^ S1817;
    assign S1819 = (X[27] & Y[1]) ^ S1818;
    assign S1820 = (X[28] & Y[0]) ^ S1819;
    assign ClmulResult[28] = S1820;
    assign S1856 = X[0] & Y[29];
    assign S1857 = (X[1] & Y[28]) ^ S1856;
    assign S1858 = (X[2] & Y[27]) ^ S1857;
    assign S1859 = (X[3] & Y[26]) ^ S1858;
    assign S1860 = (X[4] & Y[25]) ^ S1859;
    assign S1861 = (X[5] & Y[24]) ^ S1860;
    assign S1862 = (X[6] & Y[23]) ^ S1861;
    assign S1863 = (X[7] & Y[22]) ^ S1862;
    assign S1864 = (X[8] & Y[21]) ^ S1863;
    assign S1865 = (X[9] & Y[20]) ^ S1864;
    assign S1866 = (X[10] & Y[19]) ^ S1865;
    assign S1867 = (X[11] & Y[18]) ^ S1866;
    assign S1868 = (X[12] & Y[17]) ^ S1867;
    assign S1869 = (X[13] & Y[16]) ^ S1868;
    assign S1870 = (X[14] & Y[15]) ^ S1869;
    assign S1871 = (X[15] & Y[14]) ^ S1870;
    assign S1872 = (X[16] & Y[13]) ^ S1871;
    assign S1873 = (X[17] & Y[12]) ^ S1872;
    assign S1874 = (X[18] & Y[11]) ^ S1873;
    assign S1875 = (X[19] & Y[10]) ^ S1874;
    assign S1876 = (X[20] & Y[9]) ^ S1875;
    assign S1877 = (X[21] & Y[8]) ^ S1876;
    assign S1878 = (X[22] & Y[7]) ^ S1877;
    assign S1879 = (X[23] & Y[6]) ^ S1878;
    assign S1880 = (X[24] & Y[5]) ^ S1879;
    assign S1881 = (X[25] & Y[4]) ^ S1880;
    assign S1882 = (X[26] & Y[3]) ^ S1881;
    assign S1883 = (X[27] & Y[2]) ^ S1882;
    assign S1884 = (X[28] & Y[1]) ^ S1883;
    assign S1885 = (X[29] & Y[0]) ^ S1884;
    assign ClmulResult[29] = S1885;
    assign S1920 = X[0] & Y[30];
    assign S1921 = (X[1] & Y[29]) ^ S1920;
    assign S1922 = (X[2] & Y[28]) ^ S1921;
    assign S1923 = (X[3] & Y[27]) ^ S1922;
    assign S1924 = (X[4] & Y[26]) ^ S1923;
    assign S1925 = (X[5] & Y[25]) ^ S1924;
    assign S1926 = (X[6] & Y[24]) ^ S1925;
    assign S1927 = (X[7] & Y[23]) ^ S1926;
    assign S1928 = (X[8] & Y[22]) ^ S1927;
    assign S1929 = (X[9] & Y[21]) ^ S1928;
    assign S1930 = (X[10] & Y[20]) ^ S1929;
    assign S1931 = (X[11] & Y[19]) ^ S1930;
    assign S1932 = (X[12] & Y[18]) ^ S1931;
    assign S1933 = (X[13] & Y[17]) ^ S1932;
    assign S1934 = (X[14] & Y[16]) ^ S1933;
    assign S1935 = (X[15] & Y[15]) ^ S1934;
    assign S1936 = (X[16] & Y[14]) ^ S1935;
    assign S1937 = (X[17] & Y[13]) ^ S1936;
    assign S1938 = (X[18] & Y[12]) ^ S1937;
    assign S1939 = (X[19] & Y[11]) ^ S1938;
    assign S1940 = (X[20] & Y[10]) ^ S1939;
    assign S1941 = (X[21] & Y[9]) ^ S1940;
    assign S1942 = (X[22] & Y[8]) ^ S1941;
    assign S1943 = (X[23] & Y[7]) ^ S1942;
    assign S1944 = (X[24] & Y[6]) ^ S1943;
    assign S1945 = (X[25] & Y[5]) ^ S1944;
    assign S1946 = (X[26] & Y[4]) ^ S1945;
    assign S1947 = (X[27] & Y[3]) ^ S1946;
    assign S1948 = (X[28] & Y[2]) ^ S1947;
    assign S1949 = (X[29] & Y[1]) ^ S1948;
    assign S1950 = (X[30] & Y[0]) ^ S1949;
    assign ClmulResult[30] = S1950;
    assign S1984 = X[0] & Y[31];
    assign S1985 = (X[1] & Y[30]) ^ S1984;
    assign S1986 = (X[2] & Y[29]) ^ S1985;
    assign S1987 = (X[3] & Y[28]) ^ S1986;
    assign S1988 = (X[4] & Y[27]) ^ S1987;
    assign S1989 = (X[5] & Y[26]) ^ S1988;
    assign S1990 = (X[6] & Y[25]) ^ S1989;
    assign S1991 = (X[7] & Y[24]) ^ S1990;
    assign S1992 = (X[8] & Y[23]) ^ S1991;
    assign S1993 = (X[9] & Y[22]) ^ S1992;
    assign S1994 = (X[10] & Y[21]) ^ S1993;
    assign S1995 = (X[11] & Y[20]) ^ S1994;
    assign S1996 = (X[12] & Y[19]) ^ S1995;
    assign S1997 = (X[13] & Y[18]) ^ S1996;
    assign S1998 = (X[14] & Y[17]) ^ S1997;
    assign S1999 = (X[15] & Y[16]) ^ S1998;
    assign S2000 = (X[16] & Y[15]) ^ S1999;
    assign S2001 = (X[17] & Y[14]) ^ S2000;
    assign S2002 = (X[18] & Y[13]) ^ S2001;
    assign S2003 = (X[19] & Y[12]) ^ S2002;
    assign S2004 = (X[20] & Y[11]) ^ S2003;
    assign S2005 = (X[21] & Y[10]) ^ S2004;
    assign S2006 = (X[22] & Y[9]) ^ S2005;
    assign S2007 = (X[23] & Y[8]) ^ S2006;
    assign S2008 = (X[24] & Y[7]) ^ S2007;
    assign S2009 = (X[25] & Y[6]) ^ S2008;
    assign S2010 = (X[26] & Y[5]) ^ S2009;
    assign S2011 = (X[27] & Y[4]) ^ S2010;
    assign S2012 = (X[28] & Y[3]) ^ S2011;
    assign S2013 = (X[29] & Y[2]) ^ S2012;
    assign S2014 = (X[30] & Y[1]) ^ S2013;
    assign S2015 = (X[31] & Y[0]) ^ S2014;
    assign ClmulResult[31] = S2015;
    assign S2048 = X[0] & Y[32];
    assign S2049 = (X[1] & Y[31]) ^ S2048;
    assign S2050 = (X[2] & Y[30]) ^ S2049;
    assign S2051 = (X[3] & Y[29]) ^ S2050;
    assign S2052 = (X[4] & Y[28]) ^ S2051;
    assign S2053 = (X[5] & Y[27]) ^ S2052;
    assign S2054 = (X[6] & Y[26]) ^ S2053;
    assign S2055 = (X[7] & Y[25]) ^ S2054;
    assign S2056 = (X[8] & Y[24]) ^ S2055;
    assign S2057 = (X[9] & Y[23]) ^ S2056;
    assign S2058 = (X[10] & Y[22]) ^ S2057;
    assign S2059 = (X[11] & Y[21]) ^ S2058;
    assign S2060 = (X[12] & Y[20]) ^ S2059;
    assign S2061 = (X[13] & Y[19]) ^ S2060;
    assign S2062 = (X[14] & Y[18]) ^ S2061;
    assign S2063 = (X[15] & Y[17]) ^ S2062;
    assign S2064 = (X[16] & Y[16]) ^ S2063;
    assign S2065 = (X[17] & Y[15]) ^ S2064;
    assign S2066 = (X[18] & Y[14]) ^ S2065;
    assign S2067 = (X[19] & Y[13]) ^ S2066;
    assign S2068 = (X[20] & Y[12]) ^ S2067;
    assign S2069 = (X[21] & Y[11]) ^ S2068;
    assign S2070 = (X[22] & Y[10]) ^ S2069;
    assign S2071 = (X[23] & Y[9]) ^ S2070;
    assign S2072 = (X[24] & Y[8]) ^ S2071;
    assign S2073 = (X[25] & Y[7]) ^ S2072;
    assign S2074 = (X[26] & Y[6]) ^ S2073;
    assign S2075 = (X[27] & Y[5]) ^ S2074;
    assign S2076 = (X[28] & Y[4]) ^ S2075;
    assign S2077 = (X[29] & Y[3]) ^ S2076;
    assign S2078 = (X[30] & Y[2]) ^ S2077;
    assign S2079 = (X[31] & Y[1]) ^ S2078;
    assign S2080 = (X[32] & Y[0]) ^ S2079;
    assign ClmulResult[32] = S2080;
    assign S2112 = X[0] & Y[33];
    assign S2113 = (X[1] & Y[32]) ^ S2112;
    assign S2114 = (X[2] & Y[31]) ^ S2113;
    assign S2115 = (X[3] & Y[30]) ^ S2114;
    assign S2116 = (X[4] & Y[29]) ^ S2115;
    assign S2117 = (X[5] & Y[28]) ^ S2116;
    assign S2118 = (X[6] & Y[27]) ^ S2117;
    assign S2119 = (X[7] & Y[26]) ^ S2118;
    assign S2120 = (X[8] & Y[25]) ^ S2119;
    assign S2121 = (X[9] & Y[24]) ^ S2120;
    assign S2122 = (X[10] & Y[23]) ^ S2121;
    assign S2123 = (X[11] & Y[22]) ^ S2122;
    assign S2124 = (X[12] & Y[21]) ^ S2123;
    assign S2125 = (X[13] & Y[20]) ^ S2124;
    assign S2126 = (X[14] & Y[19]) ^ S2125;
    assign S2127 = (X[15] & Y[18]) ^ S2126;
    assign S2128 = (X[16] & Y[17]) ^ S2127;
    assign S2129 = (X[17] & Y[16]) ^ S2128;
    assign S2130 = (X[18] & Y[15]) ^ S2129;
    assign S2131 = (X[19] & Y[14]) ^ S2130;
    assign S2132 = (X[20] & Y[13]) ^ S2131;
    assign S2133 = (X[21] & Y[12]) ^ S2132;
    assign S2134 = (X[22] & Y[11]) ^ S2133;
    assign S2135 = (X[23] & Y[10]) ^ S2134;
    assign S2136 = (X[24] & Y[9]) ^ S2135;
    assign S2137 = (X[25] & Y[8]) ^ S2136;
    assign S2138 = (X[26] & Y[7]) ^ S2137;
    assign S2139 = (X[27] & Y[6]) ^ S2138;
    assign S2140 = (X[28] & Y[5]) ^ S2139;
    assign S2141 = (X[29] & Y[4]) ^ S2140;
    assign S2142 = (X[30] & Y[3]) ^ S2141;
    assign S2143 = (X[31] & Y[2]) ^ S2142;
    assign S2144 = (X[32] & Y[1]) ^ S2143;
    assign S2145 = (X[33] & Y[0]) ^ S2144;
    assign ClmulResult[33] = S2145;
    assign S2176 = X[0] & Y[34];
    assign S2177 = (X[1] & Y[33]) ^ S2176;
    assign S2178 = (X[2] & Y[32]) ^ S2177;
    assign S2179 = (X[3] & Y[31]) ^ S2178;
    assign S2180 = (X[4] & Y[30]) ^ S2179;
    assign S2181 = (X[5] & Y[29]) ^ S2180;
    assign S2182 = (X[6] & Y[28]) ^ S2181;
    assign S2183 = (X[7] & Y[27]) ^ S2182;
    assign S2184 = (X[8] & Y[26]) ^ S2183;
    assign S2185 = (X[9] & Y[25]) ^ S2184;
    assign S2186 = (X[10] & Y[24]) ^ S2185;
    assign S2187 = (X[11] & Y[23]) ^ S2186;
    assign S2188 = (X[12] & Y[22]) ^ S2187;
    assign S2189 = (X[13] & Y[21]) ^ S2188;
    assign S2190 = (X[14] & Y[20]) ^ S2189;
    assign S2191 = (X[15] & Y[19]) ^ S2190;
    assign S2192 = (X[16] & Y[18]) ^ S2191;
    assign S2193 = (X[17] & Y[17]) ^ S2192;
    assign S2194 = (X[18] & Y[16]) ^ S2193;
    assign S2195 = (X[19] & Y[15]) ^ S2194;
    assign S2196 = (X[20] & Y[14]) ^ S2195;
    assign S2197 = (X[21] & Y[13]) ^ S2196;
    assign S2198 = (X[22] & Y[12]) ^ S2197;
    assign S2199 = (X[23] & Y[11]) ^ S2198;
    assign S2200 = (X[24] & Y[10]) ^ S2199;
    assign S2201 = (X[25] & Y[9]) ^ S2200;
    assign S2202 = (X[26] & Y[8]) ^ S2201;
    assign S2203 = (X[27] & Y[7]) ^ S2202;
    assign S2204 = (X[28] & Y[6]) ^ S2203;
    assign S2205 = (X[29] & Y[5]) ^ S2204;
    assign S2206 = (X[30] & Y[4]) ^ S2205;
    assign S2207 = (X[31] & Y[3]) ^ S2206;
    assign S2208 = (X[32] & Y[2]) ^ S2207;
    assign S2209 = (X[33] & Y[1]) ^ S2208;
    assign S2210 = (X[34] & Y[0]) ^ S2209;
    assign ClmulResult[34] = S2210;
    assign S2240 = X[0] & Y[35];
    assign S2241 = (X[1] & Y[34]) ^ S2240;
    assign S2242 = (X[2] & Y[33]) ^ S2241;
    assign S2243 = (X[3] & Y[32]) ^ S2242;
    assign S2244 = (X[4] & Y[31]) ^ S2243;
    assign S2245 = (X[5] & Y[30]) ^ S2244;
    assign S2246 = (X[6] & Y[29]) ^ S2245;
    assign S2247 = (X[7] & Y[28]) ^ S2246;
    assign S2248 = (X[8] & Y[27]) ^ S2247;
    assign S2249 = (X[9] & Y[26]) ^ S2248;
    assign S2250 = (X[10] & Y[25]) ^ S2249;
    assign S2251 = (X[11] & Y[24]) ^ S2250;
    assign S2252 = (X[12] & Y[23]) ^ S2251;
    assign S2253 = (X[13] & Y[22]) ^ S2252;
    assign S2254 = (X[14] & Y[21]) ^ S2253;
    assign S2255 = (X[15] & Y[20]) ^ S2254;
    assign S2256 = (X[16] & Y[19]) ^ S2255;
    assign S2257 = (X[17] & Y[18]) ^ S2256;
    assign S2258 = (X[18] & Y[17]) ^ S2257;
    assign S2259 = (X[19] & Y[16]) ^ S2258;
    assign S2260 = (X[20] & Y[15]) ^ S2259;
    assign S2261 = (X[21] & Y[14]) ^ S2260;
    assign S2262 = (X[22] & Y[13]) ^ S2261;
    assign S2263 = (X[23] & Y[12]) ^ S2262;
    assign S2264 = (X[24] & Y[11]) ^ S2263;
    assign S2265 = (X[25] & Y[10]) ^ S2264;
    assign S2266 = (X[26] & Y[9]) ^ S2265;
    assign S2267 = (X[27] & Y[8]) ^ S2266;
    assign S2268 = (X[28] & Y[7]) ^ S2267;
    assign S2269 = (X[29] & Y[6]) ^ S2268;
    assign S2270 = (X[30] & Y[5]) ^ S2269;
    assign S2271 = (X[31] & Y[4]) ^ S2270;
    assign S2272 = (X[32] & Y[3]) ^ S2271;
    assign S2273 = (X[33] & Y[2]) ^ S2272;
    assign S2274 = (X[34] & Y[1]) ^ S2273;
    assign S2275 = (X[35] & Y[0]) ^ S2274;
    assign ClmulResult[35] = S2275;
    assign S2304 = X[0] & Y[36];
    assign S2305 = (X[1] & Y[35]) ^ S2304;
    assign S2306 = (X[2] & Y[34]) ^ S2305;
    assign S2307 = (X[3] & Y[33]) ^ S2306;
    assign S2308 = (X[4] & Y[32]) ^ S2307;
    assign S2309 = (X[5] & Y[31]) ^ S2308;
    assign S2310 = (X[6] & Y[30]) ^ S2309;
    assign S2311 = (X[7] & Y[29]) ^ S2310;
    assign S2312 = (X[8] & Y[28]) ^ S2311;
    assign S2313 = (X[9] & Y[27]) ^ S2312;
    assign S2314 = (X[10] & Y[26]) ^ S2313;
    assign S2315 = (X[11] & Y[25]) ^ S2314;
    assign S2316 = (X[12] & Y[24]) ^ S2315;
    assign S2317 = (X[13] & Y[23]) ^ S2316;
    assign S2318 = (X[14] & Y[22]) ^ S2317;
    assign S2319 = (X[15] & Y[21]) ^ S2318;
    assign S2320 = (X[16] & Y[20]) ^ S2319;
    assign S2321 = (X[17] & Y[19]) ^ S2320;
    assign S2322 = (X[18] & Y[18]) ^ S2321;
    assign S2323 = (X[19] & Y[17]) ^ S2322;
    assign S2324 = (X[20] & Y[16]) ^ S2323;
    assign S2325 = (X[21] & Y[15]) ^ S2324;
    assign S2326 = (X[22] & Y[14]) ^ S2325;
    assign S2327 = (X[23] & Y[13]) ^ S2326;
    assign S2328 = (X[24] & Y[12]) ^ S2327;
    assign S2329 = (X[25] & Y[11]) ^ S2328;
    assign S2330 = (X[26] & Y[10]) ^ S2329;
    assign S2331 = (X[27] & Y[9]) ^ S2330;
    assign S2332 = (X[28] & Y[8]) ^ S2331;
    assign S2333 = (X[29] & Y[7]) ^ S2332;
    assign S2334 = (X[30] & Y[6]) ^ S2333;
    assign S2335 = (X[31] & Y[5]) ^ S2334;
    assign S2336 = (X[32] & Y[4]) ^ S2335;
    assign S2337 = (X[33] & Y[3]) ^ S2336;
    assign S2338 = (X[34] & Y[2]) ^ S2337;
    assign S2339 = (X[35] & Y[1]) ^ S2338;
    assign S2340 = (X[36] & Y[0]) ^ S2339;
    assign ClmulResult[36] = S2340;
    assign S2368 = X[0] & Y[37];
    assign S2369 = (X[1] & Y[36]) ^ S2368;
    assign S2370 = (X[2] & Y[35]) ^ S2369;
    assign S2371 = (X[3] & Y[34]) ^ S2370;
    assign S2372 = (X[4] & Y[33]) ^ S2371;
    assign S2373 = (X[5] & Y[32]) ^ S2372;
    assign S2374 = (X[6] & Y[31]) ^ S2373;
    assign S2375 = (X[7] & Y[30]) ^ S2374;
    assign S2376 = (X[8] & Y[29]) ^ S2375;
    assign S2377 = (X[9] & Y[28]) ^ S2376;
    assign S2378 = (X[10] & Y[27]) ^ S2377;
    assign S2379 = (X[11] & Y[26]) ^ S2378;
    assign S2380 = (X[12] & Y[25]) ^ S2379;
    assign S2381 = (X[13] & Y[24]) ^ S2380;
    assign S2382 = (X[14] & Y[23]) ^ S2381;
    assign S2383 = (X[15] & Y[22]) ^ S2382;
    assign S2384 = (X[16] & Y[21]) ^ S2383;
    assign S2385 = (X[17] & Y[20]) ^ S2384;
    assign S2386 = (X[18] & Y[19]) ^ S2385;
    assign S2387 = (X[19] & Y[18]) ^ S2386;
    assign S2388 = (X[20] & Y[17]) ^ S2387;
    assign S2389 = (X[21] & Y[16]) ^ S2388;
    assign S2390 = (X[22] & Y[15]) ^ S2389;
    assign S2391 = (X[23] & Y[14]) ^ S2390;
    assign S2392 = (X[24] & Y[13]) ^ S2391;
    assign S2393 = (X[25] & Y[12]) ^ S2392;
    assign S2394 = (X[26] & Y[11]) ^ S2393;
    assign S2395 = (X[27] & Y[10]) ^ S2394;
    assign S2396 = (X[28] & Y[9]) ^ S2395;
    assign S2397 = (X[29] & Y[8]) ^ S2396;
    assign S2398 = (X[30] & Y[7]) ^ S2397;
    assign S2399 = (X[31] & Y[6]) ^ S2398;
    assign S2400 = (X[32] & Y[5]) ^ S2399;
    assign S2401 = (X[33] & Y[4]) ^ S2400;
    assign S2402 = (X[34] & Y[3]) ^ S2401;
    assign S2403 = (X[35] & Y[2]) ^ S2402;
    assign S2404 = (X[36] & Y[1]) ^ S2403;
    assign S2405 = (X[37] & Y[0]) ^ S2404;
    assign ClmulResult[37] = S2405;
    assign S2432 = X[0] & Y[38];
    assign S2433 = (X[1] & Y[37]) ^ S2432;
    assign S2434 = (X[2] & Y[36]) ^ S2433;
    assign S2435 = (X[3] & Y[35]) ^ S2434;
    assign S2436 = (X[4] & Y[34]) ^ S2435;
    assign S2437 = (X[5] & Y[33]) ^ S2436;
    assign S2438 = (X[6] & Y[32]) ^ S2437;
    assign S2439 = (X[7] & Y[31]) ^ S2438;
    assign S2440 = (X[8] & Y[30]) ^ S2439;
    assign S2441 = (X[9] & Y[29]) ^ S2440;
    assign S2442 = (X[10] & Y[28]) ^ S2441;
    assign S2443 = (X[11] & Y[27]) ^ S2442;
    assign S2444 = (X[12] & Y[26]) ^ S2443;
    assign S2445 = (X[13] & Y[25]) ^ S2444;
    assign S2446 = (X[14] & Y[24]) ^ S2445;
    assign S2447 = (X[15] & Y[23]) ^ S2446;
    assign S2448 = (X[16] & Y[22]) ^ S2447;
    assign S2449 = (X[17] & Y[21]) ^ S2448;
    assign S2450 = (X[18] & Y[20]) ^ S2449;
    assign S2451 = (X[19] & Y[19]) ^ S2450;
    assign S2452 = (X[20] & Y[18]) ^ S2451;
    assign S2453 = (X[21] & Y[17]) ^ S2452;
    assign S2454 = (X[22] & Y[16]) ^ S2453;
    assign S2455 = (X[23] & Y[15]) ^ S2454;
    assign S2456 = (X[24] & Y[14]) ^ S2455;
    assign S2457 = (X[25] & Y[13]) ^ S2456;
    assign S2458 = (X[26] & Y[12]) ^ S2457;
    assign S2459 = (X[27] & Y[11]) ^ S2458;
    assign S2460 = (X[28] & Y[10]) ^ S2459;
    assign S2461 = (X[29] & Y[9]) ^ S2460;
    assign S2462 = (X[30] & Y[8]) ^ S2461;
    assign S2463 = (X[31] & Y[7]) ^ S2462;
    assign S2464 = (X[32] & Y[6]) ^ S2463;
    assign S2465 = (X[33] & Y[5]) ^ S2464;
    assign S2466 = (X[34] & Y[4]) ^ S2465;
    assign S2467 = (X[35] & Y[3]) ^ S2466;
    assign S2468 = (X[36] & Y[2]) ^ S2467;
    assign S2469 = (X[37] & Y[1]) ^ S2468;
    assign S2470 = (X[38] & Y[0]) ^ S2469;
    assign ClmulResult[38] = S2470;
    assign S2496 = X[0] & Y[39];
    assign S2497 = (X[1] & Y[38]) ^ S2496;
    assign S2498 = (X[2] & Y[37]) ^ S2497;
    assign S2499 = (X[3] & Y[36]) ^ S2498;
    assign S2500 = (X[4] & Y[35]) ^ S2499;
    assign S2501 = (X[5] & Y[34]) ^ S2500;
    assign S2502 = (X[6] & Y[33]) ^ S2501;
    assign S2503 = (X[7] & Y[32]) ^ S2502;
    assign S2504 = (X[8] & Y[31]) ^ S2503;
    assign S2505 = (X[9] & Y[30]) ^ S2504;
    assign S2506 = (X[10] & Y[29]) ^ S2505;
    assign S2507 = (X[11] & Y[28]) ^ S2506;
    assign S2508 = (X[12] & Y[27]) ^ S2507;
    assign S2509 = (X[13] & Y[26]) ^ S2508;
    assign S2510 = (X[14] & Y[25]) ^ S2509;
    assign S2511 = (X[15] & Y[24]) ^ S2510;
    assign S2512 = (X[16] & Y[23]) ^ S2511;
    assign S2513 = (X[17] & Y[22]) ^ S2512;
    assign S2514 = (X[18] & Y[21]) ^ S2513;
    assign S2515 = (X[19] & Y[20]) ^ S2514;
    assign S2516 = (X[20] & Y[19]) ^ S2515;
    assign S2517 = (X[21] & Y[18]) ^ S2516;
    assign S2518 = (X[22] & Y[17]) ^ S2517;
    assign S2519 = (X[23] & Y[16]) ^ S2518;
    assign S2520 = (X[24] & Y[15]) ^ S2519;
    assign S2521 = (X[25] & Y[14]) ^ S2520;
    assign S2522 = (X[26] & Y[13]) ^ S2521;
    assign S2523 = (X[27] & Y[12]) ^ S2522;
    assign S2524 = (X[28] & Y[11]) ^ S2523;
    assign S2525 = (X[29] & Y[10]) ^ S2524;
    assign S2526 = (X[30] & Y[9]) ^ S2525;
    assign S2527 = (X[31] & Y[8]) ^ S2526;
    assign S2528 = (X[32] & Y[7]) ^ S2527;
    assign S2529 = (X[33] & Y[6]) ^ S2528;
    assign S2530 = (X[34] & Y[5]) ^ S2529;
    assign S2531 = (X[35] & Y[4]) ^ S2530;
    assign S2532 = (X[36] & Y[3]) ^ S2531;
    assign S2533 = (X[37] & Y[2]) ^ S2532;
    assign S2534 = (X[38] & Y[1]) ^ S2533;
    assign S2535 = (X[39] & Y[0]) ^ S2534;
    assign ClmulResult[39] = S2535;
    assign S2560 = X[0] & Y[40];
    assign S2561 = (X[1] & Y[39]) ^ S2560;
    assign S2562 = (X[2] & Y[38]) ^ S2561;
    assign S2563 = (X[3] & Y[37]) ^ S2562;
    assign S2564 = (X[4] & Y[36]) ^ S2563;
    assign S2565 = (X[5] & Y[35]) ^ S2564;
    assign S2566 = (X[6] & Y[34]) ^ S2565;
    assign S2567 = (X[7] & Y[33]) ^ S2566;
    assign S2568 = (X[8] & Y[32]) ^ S2567;
    assign S2569 = (X[9] & Y[31]) ^ S2568;
    assign S2570 = (X[10] & Y[30]) ^ S2569;
    assign S2571 = (X[11] & Y[29]) ^ S2570;
    assign S2572 = (X[12] & Y[28]) ^ S2571;
    assign S2573 = (X[13] & Y[27]) ^ S2572;
    assign S2574 = (X[14] & Y[26]) ^ S2573;
    assign S2575 = (X[15] & Y[25]) ^ S2574;
    assign S2576 = (X[16] & Y[24]) ^ S2575;
    assign S2577 = (X[17] & Y[23]) ^ S2576;
    assign S2578 = (X[18] & Y[22]) ^ S2577;
    assign S2579 = (X[19] & Y[21]) ^ S2578;
    assign S2580 = (X[20] & Y[20]) ^ S2579;
    assign S2581 = (X[21] & Y[19]) ^ S2580;
    assign S2582 = (X[22] & Y[18]) ^ S2581;
    assign S2583 = (X[23] & Y[17]) ^ S2582;
    assign S2584 = (X[24] & Y[16]) ^ S2583;
    assign S2585 = (X[25] & Y[15]) ^ S2584;
    assign S2586 = (X[26] & Y[14]) ^ S2585;
    assign S2587 = (X[27] & Y[13]) ^ S2586;
    assign S2588 = (X[28] & Y[12]) ^ S2587;
    assign S2589 = (X[29] & Y[11]) ^ S2588;
    assign S2590 = (X[30] & Y[10]) ^ S2589;
    assign S2591 = (X[31] & Y[9]) ^ S2590;
    assign S2592 = (X[32] & Y[8]) ^ S2591;
    assign S2593 = (X[33] & Y[7]) ^ S2592;
    assign S2594 = (X[34] & Y[6]) ^ S2593;
    assign S2595 = (X[35] & Y[5]) ^ S2594;
    assign S2596 = (X[36] & Y[4]) ^ S2595;
    assign S2597 = (X[37] & Y[3]) ^ S2596;
    assign S2598 = (X[38] & Y[2]) ^ S2597;
    assign S2599 = (X[39] & Y[1]) ^ S2598;
    assign S2600 = (X[40] & Y[0]) ^ S2599;
    assign ClmulResult[40] = S2600;
    assign S2624 = X[0] & Y[41];
    assign S2625 = (X[1] & Y[40]) ^ S2624;
    assign S2626 = (X[2] & Y[39]) ^ S2625;
    assign S2627 = (X[3] & Y[38]) ^ S2626;
    assign S2628 = (X[4] & Y[37]) ^ S2627;
    assign S2629 = (X[5] & Y[36]) ^ S2628;
    assign S2630 = (X[6] & Y[35]) ^ S2629;
    assign S2631 = (X[7] & Y[34]) ^ S2630;
    assign S2632 = (X[8] & Y[33]) ^ S2631;
    assign S2633 = (X[9] & Y[32]) ^ S2632;
    assign S2634 = (X[10] & Y[31]) ^ S2633;
    assign S2635 = (X[11] & Y[30]) ^ S2634;
    assign S2636 = (X[12] & Y[29]) ^ S2635;
    assign S2637 = (X[13] & Y[28]) ^ S2636;
    assign S2638 = (X[14] & Y[27]) ^ S2637;
    assign S2639 = (X[15] & Y[26]) ^ S2638;
    assign S2640 = (X[16] & Y[25]) ^ S2639;
    assign S2641 = (X[17] & Y[24]) ^ S2640;
    assign S2642 = (X[18] & Y[23]) ^ S2641;
    assign S2643 = (X[19] & Y[22]) ^ S2642;
    assign S2644 = (X[20] & Y[21]) ^ S2643;
    assign S2645 = (X[21] & Y[20]) ^ S2644;
    assign S2646 = (X[22] & Y[19]) ^ S2645;
    assign S2647 = (X[23] & Y[18]) ^ S2646;
    assign S2648 = (X[24] & Y[17]) ^ S2647;
    assign S2649 = (X[25] & Y[16]) ^ S2648;
    assign S2650 = (X[26] & Y[15]) ^ S2649;
    assign S2651 = (X[27] & Y[14]) ^ S2650;
    assign S2652 = (X[28] & Y[13]) ^ S2651;
    assign S2653 = (X[29] & Y[12]) ^ S2652;
    assign S2654 = (X[30] & Y[11]) ^ S2653;
    assign S2655 = (X[31] & Y[10]) ^ S2654;
    assign S2656 = (X[32] & Y[9]) ^ S2655;
    assign S2657 = (X[33] & Y[8]) ^ S2656;
    assign S2658 = (X[34] & Y[7]) ^ S2657;
    assign S2659 = (X[35] & Y[6]) ^ S2658;
    assign S2660 = (X[36] & Y[5]) ^ S2659;
    assign S2661 = (X[37] & Y[4]) ^ S2660;
    assign S2662 = (X[38] & Y[3]) ^ S2661;
    assign S2663 = (X[39] & Y[2]) ^ S2662;
    assign S2664 = (X[40] & Y[1]) ^ S2663;
    assign S2665 = (X[41] & Y[0]) ^ S2664;
    assign ClmulResult[41] = S2665;
    assign S2688 = X[0] & Y[42];
    assign S2689 = (X[1] & Y[41]) ^ S2688;
    assign S2690 = (X[2] & Y[40]) ^ S2689;
    assign S2691 = (X[3] & Y[39]) ^ S2690;
    assign S2692 = (X[4] & Y[38]) ^ S2691;
    assign S2693 = (X[5] & Y[37]) ^ S2692;
    assign S2694 = (X[6] & Y[36]) ^ S2693;
    assign S2695 = (X[7] & Y[35]) ^ S2694;
    assign S2696 = (X[8] & Y[34]) ^ S2695;
    assign S2697 = (X[9] & Y[33]) ^ S2696;
    assign S2698 = (X[10] & Y[32]) ^ S2697;
    assign S2699 = (X[11] & Y[31]) ^ S2698;
    assign S2700 = (X[12] & Y[30]) ^ S2699;
    assign S2701 = (X[13] & Y[29]) ^ S2700;
    assign S2702 = (X[14] & Y[28]) ^ S2701;
    assign S2703 = (X[15] & Y[27]) ^ S2702;
    assign S2704 = (X[16] & Y[26]) ^ S2703;
    assign S2705 = (X[17] & Y[25]) ^ S2704;
    assign S2706 = (X[18] & Y[24]) ^ S2705;
    assign S2707 = (X[19] & Y[23]) ^ S2706;
    assign S2708 = (X[20] & Y[22]) ^ S2707;
    assign S2709 = (X[21] & Y[21]) ^ S2708;
    assign S2710 = (X[22] & Y[20]) ^ S2709;
    assign S2711 = (X[23] & Y[19]) ^ S2710;
    assign S2712 = (X[24] & Y[18]) ^ S2711;
    assign S2713 = (X[25] & Y[17]) ^ S2712;
    assign S2714 = (X[26] & Y[16]) ^ S2713;
    assign S2715 = (X[27] & Y[15]) ^ S2714;
    assign S2716 = (X[28] & Y[14]) ^ S2715;
    assign S2717 = (X[29] & Y[13]) ^ S2716;
    assign S2718 = (X[30] & Y[12]) ^ S2717;
    assign S2719 = (X[31] & Y[11]) ^ S2718;
    assign S2720 = (X[32] & Y[10]) ^ S2719;
    assign S2721 = (X[33] & Y[9]) ^ S2720;
    assign S2722 = (X[34] & Y[8]) ^ S2721;
    assign S2723 = (X[35] & Y[7]) ^ S2722;
    assign S2724 = (X[36] & Y[6]) ^ S2723;
    assign S2725 = (X[37] & Y[5]) ^ S2724;
    assign S2726 = (X[38] & Y[4]) ^ S2725;
    assign S2727 = (X[39] & Y[3]) ^ S2726;
    assign S2728 = (X[40] & Y[2]) ^ S2727;
    assign S2729 = (X[41] & Y[1]) ^ S2728;
    assign S2730 = (X[42] & Y[0]) ^ S2729;
    assign ClmulResult[42] = S2730;
    assign S2752 = X[0] & Y[43];
    assign S2753 = (X[1] & Y[42]) ^ S2752;
    assign S2754 = (X[2] & Y[41]) ^ S2753;
    assign S2755 = (X[3] & Y[40]) ^ S2754;
    assign S2756 = (X[4] & Y[39]) ^ S2755;
    assign S2757 = (X[5] & Y[38]) ^ S2756;
    assign S2758 = (X[6] & Y[37]) ^ S2757;
    assign S2759 = (X[7] & Y[36]) ^ S2758;
    assign S2760 = (X[8] & Y[35]) ^ S2759;
    assign S2761 = (X[9] & Y[34]) ^ S2760;
    assign S2762 = (X[10] & Y[33]) ^ S2761;
    assign S2763 = (X[11] & Y[32]) ^ S2762;
    assign S2764 = (X[12] & Y[31]) ^ S2763;
    assign S2765 = (X[13] & Y[30]) ^ S2764;
    assign S2766 = (X[14] & Y[29]) ^ S2765;
    assign S2767 = (X[15] & Y[28]) ^ S2766;
    assign S2768 = (X[16] & Y[27]) ^ S2767;
    assign S2769 = (X[17] & Y[26]) ^ S2768;
    assign S2770 = (X[18] & Y[25]) ^ S2769;
    assign S2771 = (X[19] & Y[24]) ^ S2770;
    assign S2772 = (X[20] & Y[23]) ^ S2771;
    assign S2773 = (X[21] & Y[22]) ^ S2772;
    assign S2774 = (X[22] & Y[21]) ^ S2773;
    assign S2775 = (X[23] & Y[20]) ^ S2774;
    assign S2776 = (X[24] & Y[19]) ^ S2775;
    assign S2777 = (X[25] & Y[18]) ^ S2776;
    assign S2778 = (X[26] & Y[17]) ^ S2777;
    assign S2779 = (X[27] & Y[16]) ^ S2778;
    assign S2780 = (X[28] & Y[15]) ^ S2779;
    assign S2781 = (X[29] & Y[14]) ^ S2780;
    assign S2782 = (X[30] & Y[13]) ^ S2781;
    assign S2783 = (X[31] & Y[12]) ^ S2782;
    assign S2784 = (X[32] & Y[11]) ^ S2783;
    assign S2785 = (X[33] & Y[10]) ^ S2784;
    assign S2786 = (X[34] & Y[9]) ^ S2785;
    assign S2787 = (X[35] & Y[8]) ^ S2786;
    assign S2788 = (X[36] & Y[7]) ^ S2787;
    assign S2789 = (X[37] & Y[6]) ^ S2788;
    assign S2790 = (X[38] & Y[5]) ^ S2789;
    assign S2791 = (X[39] & Y[4]) ^ S2790;
    assign S2792 = (X[40] & Y[3]) ^ S2791;
    assign S2793 = (X[41] & Y[2]) ^ S2792;
    assign S2794 = (X[42] & Y[1]) ^ S2793;
    assign S2795 = (X[43] & Y[0]) ^ S2794;
    assign ClmulResult[43] = S2795;
    assign S2816 = X[0] & Y[44];
    assign S2817 = (X[1] & Y[43]) ^ S2816;
    assign S2818 = (X[2] & Y[42]) ^ S2817;
    assign S2819 = (X[3] & Y[41]) ^ S2818;
    assign S2820 = (X[4] & Y[40]) ^ S2819;
    assign S2821 = (X[5] & Y[39]) ^ S2820;
    assign S2822 = (X[6] & Y[38]) ^ S2821;
    assign S2823 = (X[7] & Y[37]) ^ S2822;
    assign S2824 = (X[8] & Y[36]) ^ S2823;
    assign S2825 = (X[9] & Y[35]) ^ S2824;
    assign S2826 = (X[10] & Y[34]) ^ S2825;
    assign S2827 = (X[11] & Y[33]) ^ S2826;
    assign S2828 = (X[12] & Y[32]) ^ S2827;
    assign S2829 = (X[13] & Y[31]) ^ S2828;
    assign S2830 = (X[14] & Y[30]) ^ S2829;
    assign S2831 = (X[15] & Y[29]) ^ S2830;
    assign S2832 = (X[16] & Y[28]) ^ S2831;
    assign S2833 = (X[17] & Y[27]) ^ S2832;
    assign S2834 = (X[18] & Y[26]) ^ S2833;
    assign S2835 = (X[19] & Y[25]) ^ S2834;
    assign S2836 = (X[20] & Y[24]) ^ S2835;
    assign S2837 = (X[21] & Y[23]) ^ S2836;
    assign S2838 = (X[22] & Y[22]) ^ S2837;
    assign S2839 = (X[23] & Y[21]) ^ S2838;
    assign S2840 = (X[24] & Y[20]) ^ S2839;
    assign S2841 = (X[25] & Y[19]) ^ S2840;
    assign S2842 = (X[26] & Y[18]) ^ S2841;
    assign S2843 = (X[27] & Y[17]) ^ S2842;
    assign S2844 = (X[28] & Y[16]) ^ S2843;
    assign S2845 = (X[29] & Y[15]) ^ S2844;
    assign S2846 = (X[30] & Y[14]) ^ S2845;
    assign S2847 = (X[31] & Y[13]) ^ S2846;
    assign S2848 = (X[32] & Y[12]) ^ S2847;
    assign S2849 = (X[33] & Y[11]) ^ S2848;
    assign S2850 = (X[34] & Y[10]) ^ S2849;
    assign S2851 = (X[35] & Y[9]) ^ S2850;
    assign S2852 = (X[36] & Y[8]) ^ S2851;
    assign S2853 = (X[37] & Y[7]) ^ S2852;
    assign S2854 = (X[38] & Y[6]) ^ S2853;
    assign S2855 = (X[39] & Y[5]) ^ S2854;
    assign S2856 = (X[40] & Y[4]) ^ S2855;
    assign S2857 = (X[41] & Y[3]) ^ S2856;
    assign S2858 = (X[42] & Y[2]) ^ S2857;
    assign S2859 = (X[43] & Y[1]) ^ S2858;
    assign S2860 = (X[44] & Y[0]) ^ S2859;
    assign ClmulResult[44] = S2860;
    assign S2880 = X[0] & Y[45];
    assign S2881 = (X[1] & Y[44]) ^ S2880;
    assign S2882 = (X[2] & Y[43]) ^ S2881;
    assign S2883 = (X[3] & Y[42]) ^ S2882;
    assign S2884 = (X[4] & Y[41]) ^ S2883;
    assign S2885 = (X[5] & Y[40]) ^ S2884;
    assign S2886 = (X[6] & Y[39]) ^ S2885;
    assign S2887 = (X[7] & Y[38]) ^ S2886;
    assign S2888 = (X[8] & Y[37]) ^ S2887;
    assign S2889 = (X[9] & Y[36]) ^ S2888;
    assign S2890 = (X[10] & Y[35]) ^ S2889;
    assign S2891 = (X[11] & Y[34]) ^ S2890;
    assign S2892 = (X[12] & Y[33]) ^ S2891;
    assign S2893 = (X[13] & Y[32]) ^ S2892;
    assign S2894 = (X[14] & Y[31]) ^ S2893;
    assign S2895 = (X[15] & Y[30]) ^ S2894;
    assign S2896 = (X[16] & Y[29]) ^ S2895;
    assign S2897 = (X[17] & Y[28]) ^ S2896;
    assign S2898 = (X[18] & Y[27]) ^ S2897;
    assign S2899 = (X[19] & Y[26]) ^ S2898;
    assign S2900 = (X[20] & Y[25]) ^ S2899;
    assign S2901 = (X[21] & Y[24]) ^ S2900;
    assign S2902 = (X[22] & Y[23]) ^ S2901;
    assign S2903 = (X[23] & Y[22]) ^ S2902;
    assign S2904 = (X[24] & Y[21]) ^ S2903;
    assign S2905 = (X[25] & Y[20]) ^ S2904;
    assign S2906 = (X[26] & Y[19]) ^ S2905;
    assign S2907 = (X[27] & Y[18]) ^ S2906;
    assign S2908 = (X[28] & Y[17]) ^ S2907;
    assign S2909 = (X[29] & Y[16]) ^ S2908;
    assign S2910 = (X[30] & Y[15]) ^ S2909;
    assign S2911 = (X[31] & Y[14]) ^ S2910;
    assign S2912 = (X[32] & Y[13]) ^ S2911;
    assign S2913 = (X[33] & Y[12]) ^ S2912;
    assign S2914 = (X[34] & Y[11]) ^ S2913;
    assign S2915 = (X[35] & Y[10]) ^ S2914;
    assign S2916 = (X[36] & Y[9]) ^ S2915;
    assign S2917 = (X[37] & Y[8]) ^ S2916;
    assign S2918 = (X[38] & Y[7]) ^ S2917;
    assign S2919 = (X[39] & Y[6]) ^ S2918;
    assign S2920 = (X[40] & Y[5]) ^ S2919;
    assign S2921 = (X[41] & Y[4]) ^ S2920;
    assign S2922 = (X[42] & Y[3]) ^ S2921;
    assign S2923 = (X[43] & Y[2]) ^ S2922;
    assign S2924 = (X[44] & Y[1]) ^ S2923;
    assign S2925 = (X[45] & Y[0]) ^ S2924;
    assign ClmulResult[45] = S2925;
    assign S2944 = X[0] & Y[46];
    assign S2945 = (X[1] & Y[45]) ^ S2944;
    assign S2946 = (X[2] & Y[44]) ^ S2945;
    assign S2947 = (X[3] & Y[43]) ^ S2946;
    assign S2948 = (X[4] & Y[42]) ^ S2947;
    assign S2949 = (X[5] & Y[41]) ^ S2948;
    assign S2950 = (X[6] & Y[40]) ^ S2949;
    assign S2951 = (X[7] & Y[39]) ^ S2950;
    assign S2952 = (X[8] & Y[38]) ^ S2951;
    assign S2953 = (X[9] & Y[37]) ^ S2952;
    assign S2954 = (X[10] & Y[36]) ^ S2953;
    assign S2955 = (X[11] & Y[35]) ^ S2954;
    assign S2956 = (X[12] & Y[34]) ^ S2955;
    assign S2957 = (X[13] & Y[33]) ^ S2956;
    assign S2958 = (X[14] & Y[32]) ^ S2957;
    assign S2959 = (X[15] & Y[31]) ^ S2958;
    assign S2960 = (X[16] & Y[30]) ^ S2959;
    assign S2961 = (X[17] & Y[29]) ^ S2960;
    assign S2962 = (X[18] & Y[28]) ^ S2961;
    assign S2963 = (X[19] & Y[27]) ^ S2962;
    assign S2964 = (X[20] & Y[26]) ^ S2963;
    assign S2965 = (X[21] & Y[25]) ^ S2964;
    assign S2966 = (X[22] & Y[24]) ^ S2965;
    assign S2967 = (X[23] & Y[23]) ^ S2966;
    assign S2968 = (X[24] & Y[22]) ^ S2967;
    assign S2969 = (X[25] & Y[21]) ^ S2968;
    assign S2970 = (X[26] & Y[20]) ^ S2969;
    assign S2971 = (X[27] & Y[19]) ^ S2970;
    assign S2972 = (X[28] & Y[18]) ^ S2971;
    assign S2973 = (X[29] & Y[17]) ^ S2972;
    assign S2974 = (X[30] & Y[16]) ^ S2973;
    assign S2975 = (X[31] & Y[15]) ^ S2974;
    assign S2976 = (X[32] & Y[14]) ^ S2975;
    assign S2977 = (X[33] & Y[13]) ^ S2976;
    assign S2978 = (X[34] & Y[12]) ^ S2977;
    assign S2979 = (X[35] & Y[11]) ^ S2978;
    assign S2980 = (X[36] & Y[10]) ^ S2979;
    assign S2981 = (X[37] & Y[9]) ^ S2980;
    assign S2982 = (X[38] & Y[8]) ^ S2981;
    assign S2983 = (X[39] & Y[7]) ^ S2982;
    assign S2984 = (X[40] & Y[6]) ^ S2983;
    assign S2985 = (X[41] & Y[5]) ^ S2984;
    assign S2986 = (X[42] & Y[4]) ^ S2985;
    assign S2987 = (X[43] & Y[3]) ^ S2986;
    assign S2988 = (X[44] & Y[2]) ^ S2987;
    assign S2989 = (X[45] & Y[1]) ^ S2988;
    assign S2990 = (X[46] & Y[0]) ^ S2989;
    assign ClmulResult[46] = S2990;
    assign S3008 = X[0] & Y[47];
    assign S3009 = (X[1] & Y[46]) ^ S3008;
    assign S3010 = (X[2] & Y[45]) ^ S3009;
    assign S3011 = (X[3] & Y[44]) ^ S3010;
    assign S3012 = (X[4] & Y[43]) ^ S3011;
    assign S3013 = (X[5] & Y[42]) ^ S3012;
    assign S3014 = (X[6] & Y[41]) ^ S3013;
    assign S3015 = (X[7] & Y[40]) ^ S3014;
    assign S3016 = (X[8] & Y[39]) ^ S3015;
    assign S3017 = (X[9] & Y[38]) ^ S3016;
    assign S3018 = (X[10] & Y[37]) ^ S3017;
    assign S3019 = (X[11] & Y[36]) ^ S3018;
    assign S3020 = (X[12] & Y[35]) ^ S3019;
    assign S3021 = (X[13] & Y[34]) ^ S3020;
    assign S3022 = (X[14] & Y[33]) ^ S3021;
    assign S3023 = (X[15] & Y[32]) ^ S3022;
    assign S3024 = (X[16] & Y[31]) ^ S3023;
    assign S3025 = (X[17] & Y[30]) ^ S3024;
    assign S3026 = (X[18] & Y[29]) ^ S3025;
    assign S3027 = (X[19] & Y[28]) ^ S3026;
    assign S3028 = (X[20] & Y[27]) ^ S3027;
    assign S3029 = (X[21] & Y[26]) ^ S3028;
    assign S3030 = (X[22] & Y[25]) ^ S3029;
    assign S3031 = (X[23] & Y[24]) ^ S3030;
    assign S3032 = (X[24] & Y[23]) ^ S3031;
    assign S3033 = (X[25] & Y[22]) ^ S3032;
    assign S3034 = (X[26] & Y[21]) ^ S3033;
    assign S3035 = (X[27] & Y[20]) ^ S3034;
    assign S3036 = (X[28] & Y[19]) ^ S3035;
    assign S3037 = (X[29] & Y[18]) ^ S3036;
    assign S3038 = (X[30] & Y[17]) ^ S3037;
    assign S3039 = (X[31] & Y[16]) ^ S3038;
    assign S3040 = (X[32] & Y[15]) ^ S3039;
    assign S3041 = (X[33] & Y[14]) ^ S3040;
    assign S3042 = (X[34] & Y[13]) ^ S3041;
    assign S3043 = (X[35] & Y[12]) ^ S3042;
    assign S3044 = (X[36] & Y[11]) ^ S3043;
    assign S3045 = (X[37] & Y[10]) ^ S3044;
    assign S3046 = (X[38] & Y[9]) ^ S3045;
    assign S3047 = (X[39] & Y[8]) ^ S3046;
    assign S3048 = (X[40] & Y[7]) ^ S3047;
    assign S3049 = (X[41] & Y[6]) ^ S3048;
    assign S3050 = (X[42] & Y[5]) ^ S3049;
    assign S3051 = (X[43] & Y[4]) ^ S3050;
    assign S3052 = (X[44] & Y[3]) ^ S3051;
    assign S3053 = (X[45] & Y[2]) ^ S3052;
    assign S3054 = (X[46] & Y[1]) ^ S3053;
    assign S3055 = (X[47] & Y[0]) ^ S3054;
    assign ClmulResult[47] = S3055;
    assign S3072 = X[0] & Y[48];
    assign S3073 = (X[1] & Y[47]) ^ S3072;
    assign S3074 = (X[2] & Y[46]) ^ S3073;
    assign S3075 = (X[3] & Y[45]) ^ S3074;
    assign S3076 = (X[4] & Y[44]) ^ S3075;
    assign S3077 = (X[5] & Y[43]) ^ S3076;
    assign S3078 = (X[6] & Y[42]) ^ S3077;
    assign S3079 = (X[7] & Y[41]) ^ S3078;
    assign S3080 = (X[8] & Y[40]) ^ S3079;
    assign S3081 = (X[9] & Y[39]) ^ S3080;
    assign S3082 = (X[10] & Y[38]) ^ S3081;
    assign S3083 = (X[11] & Y[37]) ^ S3082;
    assign S3084 = (X[12] & Y[36]) ^ S3083;
    assign S3085 = (X[13] & Y[35]) ^ S3084;
    assign S3086 = (X[14] & Y[34]) ^ S3085;
    assign S3087 = (X[15] & Y[33]) ^ S3086;
    assign S3088 = (X[16] & Y[32]) ^ S3087;
    assign S3089 = (X[17] & Y[31]) ^ S3088;
    assign S3090 = (X[18] & Y[30]) ^ S3089;
    assign S3091 = (X[19] & Y[29]) ^ S3090;
    assign S3092 = (X[20] & Y[28]) ^ S3091;
    assign S3093 = (X[21] & Y[27]) ^ S3092;
    assign S3094 = (X[22] & Y[26]) ^ S3093;
    assign S3095 = (X[23] & Y[25]) ^ S3094;
    assign S3096 = (X[24] & Y[24]) ^ S3095;
    assign S3097 = (X[25] & Y[23]) ^ S3096;
    assign S3098 = (X[26] & Y[22]) ^ S3097;
    assign S3099 = (X[27] & Y[21]) ^ S3098;
    assign S3100 = (X[28] & Y[20]) ^ S3099;
    assign S3101 = (X[29] & Y[19]) ^ S3100;
    assign S3102 = (X[30] & Y[18]) ^ S3101;
    assign S3103 = (X[31] & Y[17]) ^ S3102;
    assign S3104 = (X[32] & Y[16]) ^ S3103;
    assign S3105 = (X[33] & Y[15]) ^ S3104;
    assign S3106 = (X[34] & Y[14]) ^ S3105;
    assign S3107 = (X[35] & Y[13]) ^ S3106;
    assign S3108 = (X[36] & Y[12]) ^ S3107;
    assign S3109 = (X[37] & Y[11]) ^ S3108;
    assign S3110 = (X[38] & Y[10]) ^ S3109;
    assign S3111 = (X[39] & Y[9]) ^ S3110;
    assign S3112 = (X[40] & Y[8]) ^ S3111;
    assign S3113 = (X[41] & Y[7]) ^ S3112;
    assign S3114 = (X[42] & Y[6]) ^ S3113;
    assign S3115 = (X[43] & Y[5]) ^ S3114;
    assign S3116 = (X[44] & Y[4]) ^ S3115;
    assign S3117 = (X[45] & Y[3]) ^ S3116;
    assign S3118 = (X[46] & Y[2]) ^ S3117;
    assign S3119 = (X[47] & Y[1]) ^ S3118;
    assign S3120 = (X[48] & Y[0]) ^ S3119;
    assign ClmulResult[48] = S3120;
    assign S3136 = X[0] & Y[49];
    assign S3137 = (X[1] & Y[48]) ^ S3136;
    assign S3138 = (X[2] & Y[47]) ^ S3137;
    assign S3139 = (X[3] & Y[46]) ^ S3138;
    assign S3140 = (X[4] & Y[45]) ^ S3139;
    assign S3141 = (X[5] & Y[44]) ^ S3140;
    assign S3142 = (X[6] & Y[43]) ^ S3141;
    assign S3143 = (X[7] & Y[42]) ^ S3142;
    assign S3144 = (X[8] & Y[41]) ^ S3143;
    assign S3145 = (X[9] & Y[40]) ^ S3144;
    assign S3146 = (X[10] & Y[39]) ^ S3145;
    assign S3147 = (X[11] & Y[38]) ^ S3146;
    assign S3148 = (X[12] & Y[37]) ^ S3147;
    assign S3149 = (X[13] & Y[36]) ^ S3148;
    assign S3150 = (X[14] & Y[35]) ^ S3149;
    assign S3151 = (X[15] & Y[34]) ^ S3150;
    assign S3152 = (X[16] & Y[33]) ^ S3151;
    assign S3153 = (X[17] & Y[32]) ^ S3152;
    assign S3154 = (X[18] & Y[31]) ^ S3153;
    assign S3155 = (X[19] & Y[30]) ^ S3154;
    assign S3156 = (X[20] & Y[29]) ^ S3155;
    assign S3157 = (X[21] & Y[28]) ^ S3156;
    assign S3158 = (X[22] & Y[27]) ^ S3157;
    assign S3159 = (X[23] & Y[26]) ^ S3158;
    assign S3160 = (X[24] & Y[25]) ^ S3159;
    assign S3161 = (X[25] & Y[24]) ^ S3160;
    assign S3162 = (X[26] & Y[23]) ^ S3161;
    assign S3163 = (X[27] & Y[22]) ^ S3162;
    assign S3164 = (X[28] & Y[21]) ^ S3163;
    assign S3165 = (X[29] & Y[20]) ^ S3164;
    assign S3166 = (X[30] & Y[19]) ^ S3165;
    assign S3167 = (X[31] & Y[18]) ^ S3166;
    assign S3168 = (X[32] & Y[17]) ^ S3167;
    assign S3169 = (X[33] & Y[16]) ^ S3168;
    assign S3170 = (X[34] & Y[15]) ^ S3169;
    assign S3171 = (X[35] & Y[14]) ^ S3170;
    assign S3172 = (X[36] & Y[13]) ^ S3171;
    assign S3173 = (X[37] & Y[12]) ^ S3172;
    assign S3174 = (X[38] & Y[11]) ^ S3173;
    assign S3175 = (X[39] & Y[10]) ^ S3174;
    assign S3176 = (X[40] & Y[9]) ^ S3175;
    assign S3177 = (X[41] & Y[8]) ^ S3176;
    assign S3178 = (X[42] & Y[7]) ^ S3177;
    assign S3179 = (X[43] & Y[6]) ^ S3178;
    assign S3180 = (X[44] & Y[5]) ^ S3179;
    assign S3181 = (X[45] & Y[4]) ^ S3180;
    assign S3182 = (X[46] & Y[3]) ^ S3181;
    assign S3183 = (X[47] & Y[2]) ^ S3182;
    assign S3184 = (X[48] & Y[1]) ^ S3183;
    assign S3185 = (X[49] & Y[0]) ^ S3184;
    assign ClmulResult[49] = S3185;
    assign S3200 = X[0] & Y[50];
    assign S3201 = (X[1] & Y[49]) ^ S3200;
    assign S3202 = (X[2] & Y[48]) ^ S3201;
    assign S3203 = (X[3] & Y[47]) ^ S3202;
    assign S3204 = (X[4] & Y[46]) ^ S3203;
    assign S3205 = (X[5] & Y[45]) ^ S3204;
    assign S3206 = (X[6] & Y[44]) ^ S3205;
    assign S3207 = (X[7] & Y[43]) ^ S3206;
    assign S3208 = (X[8] & Y[42]) ^ S3207;
    assign S3209 = (X[9] & Y[41]) ^ S3208;
    assign S3210 = (X[10] & Y[40]) ^ S3209;
    assign S3211 = (X[11] & Y[39]) ^ S3210;
    assign S3212 = (X[12] & Y[38]) ^ S3211;
    assign S3213 = (X[13] & Y[37]) ^ S3212;
    assign S3214 = (X[14] & Y[36]) ^ S3213;
    assign S3215 = (X[15] & Y[35]) ^ S3214;
    assign S3216 = (X[16] & Y[34]) ^ S3215;
    assign S3217 = (X[17] & Y[33]) ^ S3216;
    assign S3218 = (X[18] & Y[32]) ^ S3217;
    assign S3219 = (X[19] & Y[31]) ^ S3218;
    assign S3220 = (X[20] & Y[30]) ^ S3219;
    assign S3221 = (X[21] & Y[29]) ^ S3220;
    assign S3222 = (X[22] & Y[28]) ^ S3221;
    assign S3223 = (X[23] & Y[27]) ^ S3222;
    assign S3224 = (X[24] & Y[26]) ^ S3223;
    assign S3225 = (X[25] & Y[25]) ^ S3224;
    assign S3226 = (X[26] & Y[24]) ^ S3225;
    assign S3227 = (X[27] & Y[23]) ^ S3226;
    assign S3228 = (X[28] & Y[22]) ^ S3227;
    assign S3229 = (X[29] & Y[21]) ^ S3228;
    assign S3230 = (X[30] & Y[20]) ^ S3229;
    assign S3231 = (X[31] & Y[19]) ^ S3230;
    assign S3232 = (X[32] & Y[18]) ^ S3231;
    assign S3233 = (X[33] & Y[17]) ^ S3232;
    assign S3234 = (X[34] & Y[16]) ^ S3233;
    assign S3235 = (X[35] & Y[15]) ^ S3234;
    assign S3236 = (X[36] & Y[14]) ^ S3235;
    assign S3237 = (X[37] & Y[13]) ^ S3236;
    assign S3238 = (X[38] & Y[12]) ^ S3237;
    assign S3239 = (X[39] & Y[11]) ^ S3238;
    assign S3240 = (X[40] & Y[10]) ^ S3239;
    assign S3241 = (X[41] & Y[9]) ^ S3240;
    assign S3242 = (X[42] & Y[8]) ^ S3241;
    assign S3243 = (X[43] & Y[7]) ^ S3242;
    assign S3244 = (X[44] & Y[6]) ^ S3243;
    assign S3245 = (X[45] & Y[5]) ^ S3244;
    assign S3246 = (X[46] & Y[4]) ^ S3245;
    assign S3247 = (X[47] & Y[3]) ^ S3246;
    assign S3248 = (X[48] & Y[2]) ^ S3247;
    assign S3249 = (X[49] & Y[1]) ^ S3248;
    assign S3250 = (X[50] & Y[0]) ^ S3249;
    assign ClmulResult[50] = S3250;
    assign S3264 = X[0] & Y[51];
    assign S3265 = (X[1] & Y[50]) ^ S3264;
    assign S3266 = (X[2] & Y[49]) ^ S3265;
    assign S3267 = (X[3] & Y[48]) ^ S3266;
    assign S3268 = (X[4] & Y[47]) ^ S3267;
    assign S3269 = (X[5] & Y[46]) ^ S3268;
    assign S3270 = (X[6] & Y[45]) ^ S3269;
    assign S3271 = (X[7] & Y[44]) ^ S3270;
    assign S3272 = (X[8] & Y[43]) ^ S3271;
    assign S3273 = (X[9] & Y[42]) ^ S3272;
    assign S3274 = (X[10] & Y[41]) ^ S3273;
    assign S3275 = (X[11] & Y[40]) ^ S3274;
    assign S3276 = (X[12] & Y[39]) ^ S3275;
    assign S3277 = (X[13] & Y[38]) ^ S3276;
    assign S3278 = (X[14] & Y[37]) ^ S3277;
    assign S3279 = (X[15] & Y[36]) ^ S3278;
    assign S3280 = (X[16] & Y[35]) ^ S3279;
    assign S3281 = (X[17] & Y[34]) ^ S3280;
    assign S3282 = (X[18] & Y[33]) ^ S3281;
    assign S3283 = (X[19] & Y[32]) ^ S3282;
    assign S3284 = (X[20] & Y[31]) ^ S3283;
    assign S3285 = (X[21] & Y[30]) ^ S3284;
    assign S3286 = (X[22] & Y[29]) ^ S3285;
    assign S3287 = (X[23] & Y[28]) ^ S3286;
    assign S3288 = (X[24] & Y[27]) ^ S3287;
    assign S3289 = (X[25] & Y[26]) ^ S3288;
    assign S3290 = (X[26] & Y[25]) ^ S3289;
    assign S3291 = (X[27] & Y[24]) ^ S3290;
    assign S3292 = (X[28] & Y[23]) ^ S3291;
    assign S3293 = (X[29] & Y[22]) ^ S3292;
    assign S3294 = (X[30] & Y[21]) ^ S3293;
    assign S3295 = (X[31] & Y[20]) ^ S3294;
    assign S3296 = (X[32] & Y[19]) ^ S3295;
    assign S3297 = (X[33] & Y[18]) ^ S3296;
    assign S3298 = (X[34] & Y[17]) ^ S3297;
    assign S3299 = (X[35] & Y[16]) ^ S3298;
    assign S3300 = (X[36] & Y[15]) ^ S3299;
    assign S3301 = (X[37] & Y[14]) ^ S3300;
    assign S3302 = (X[38] & Y[13]) ^ S3301;
    assign S3303 = (X[39] & Y[12]) ^ S3302;
    assign S3304 = (X[40] & Y[11]) ^ S3303;
    assign S3305 = (X[41] & Y[10]) ^ S3304;
    assign S3306 = (X[42] & Y[9]) ^ S3305;
    assign S3307 = (X[43] & Y[8]) ^ S3306;
    assign S3308 = (X[44] & Y[7]) ^ S3307;
    assign S3309 = (X[45] & Y[6]) ^ S3308;
    assign S3310 = (X[46] & Y[5]) ^ S3309;
    assign S3311 = (X[47] & Y[4]) ^ S3310;
    assign S3312 = (X[48] & Y[3]) ^ S3311;
    assign S3313 = (X[49] & Y[2]) ^ S3312;
    assign S3314 = (X[50] & Y[1]) ^ S3313;
    assign S3315 = (X[51] & Y[0]) ^ S3314;
    assign ClmulResult[51] = S3315;
    assign S3328 = X[0] & Y[52];
    assign S3329 = (X[1] & Y[51]) ^ S3328;
    assign S3330 = (X[2] & Y[50]) ^ S3329;
    assign S3331 = (X[3] & Y[49]) ^ S3330;
    assign S3332 = (X[4] & Y[48]) ^ S3331;
    assign S3333 = (X[5] & Y[47]) ^ S3332;
    assign S3334 = (X[6] & Y[46]) ^ S3333;
    assign S3335 = (X[7] & Y[45]) ^ S3334;
    assign S3336 = (X[8] & Y[44]) ^ S3335;
    assign S3337 = (X[9] & Y[43]) ^ S3336;
    assign S3338 = (X[10] & Y[42]) ^ S3337;
    assign S3339 = (X[11] & Y[41]) ^ S3338;
    assign S3340 = (X[12] & Y[40]) ^ S3339;
    assign S3341 = (X[13] & Y[39]) ^ S3340;
    assign S3342 = (X[14] & Y[38]) ^ S3341;
    assign S3343 = (X[15] & Y[37]) ^ S3342;
    assign S3344 = (X[16] & Y[36]) ^ S3343;
    assign S3345 = (X[17] & Y[35]) ^ S3344;
    assign S3346 = (X[18] & Y[34]) ^ S3345;
    assign S3347 = (X[19] & Y[33]) ^ S3346;
    assign S3348 = (X[20] & Y[32]) ^ S3347;
    assign S3349 = (X[21] & Y[31]) ^ S3348;
    assign S3350 = (X[22] & Y[30]) ^ S3349;
    assign S3351 = (X[23] & Y[29]) ^ S3350;
    assign S3352 = (X[24] & Y[28]) ^ S3351;
    assign S3353 = (X[25] & Y[27]) ^ S3352;
    assign S3354 = (X[26] & Y[26]) ^ S3353;
    assign S3355 = (X[27] & Y[25]) ^ S3354;
    assign S3356 = (X[28] & Y[24]) ^ S3355;
    assign S3357 = (X[29] & Y[23]) ^ S3356;
    assign S3358 = (X[30] & Y[22]) ^ S3357;
    assign S3359 = (X[31] & Y[21]) ^ S3358;
    assign S3360 = (X[32] & Y[20]) ^ S3359;
    assign S3361 = (X[33] & Y[19]) ^ S3360;
    assign S3362 = (X[34] & Y[18]) ^ S3361;
    assign S3363 = (X[35] & Y[17]) ^ S3362;
    assign S3364 = (X[36] & Y[16]) ^ S3363;
    assign S3365 = (X[37] & Y[15]) ^ S3364;
    assign S3366 = (X[38] & Y[14]) ^ S3365;
    assign S3367 = (X[39] & Y[13]) ^ S3366;
    assign S3368 = (X[40] & Y[12]) ^ S3367;
    assign S3369 = (X[41] & Y[11]) ^ S3368;
    assign S3370 = (X[42] & Y[10]) ^ S3369;
    assign S3371 = (X[43] & Y[9]) ^ S3370;
    assign S3372 = (X[44] & Y[8]) ^ S3371;
    assign S3373 = (X[45] & Y[7]) ^ S3372;
    assign S3374 = (X[46] & Y[6]) ^ S3373;
    assign S3375 = (X[47] & Y[5]) ^ S3374;
    assign S3376 = (X[48] & Y[4]) ^ S3375;
    assign S3377 = (X[49] & Y[3]) ^ S3376;
    assign S3378 = (X[50] & Y[2]) ^ S3377;
    assign S3379 = (X[51] & Y[1]) ^ S3378;
    assign S3380 = (X[52] & Y[0]) ^ S3379;
    assign ClmulResult[52] = S3380;
    assign S3392 = X[0] & Y[53];
    assign S3393 = (X[1] & Y[52]) ^ S3392;
    assign S3394 = (X[2] & Y[51]) ^ S3393;
    assign S3395 = (X[3] & Y[50]) ^ S3394;
    assign S3396 = (X[4] & Y[49]) ^ S3395;
    assign S3397 = (X[5] & Y[48]) ^ S3396;
    assign S3398 = (X[6] & Y[47]) ^ S3397;
    assign S3399 = (X[7] & Y[46]) ^ S3398;
    assign S3400 = (X[8] & Y[45]) ^ S3399;
    assign S3401 = (X[9] & Y[44]) ^ S3400;
    assign S3402 = (X[10] & Y[43]) ^ S3401;
    assign S3403 = (X[11] & Y[42]) ^ S3402;
    assign S3404 = (X[12] & Y[41]) ^ S3403;
    assign S3405 = (X[13] & Y[40]) ^ S3404;
    assign S3406 = (X[14] & Y[39]) ^ S3405;
    assign S3407 = (X[15] & Y[38]) ^ S3406;
    assign S3408 = (X[16] & Y[37]) ^ S3407;
    assign S3409 = (X[17] & Y[36]) ^ S3408;
    assign S3410 = (X[18] & Y[35]) ^ S3409;
    assign S3411 = (X[19] & Y[34]) ^ S3410;
    assign S3412 = (X[20] & Y[33]) ^ S3411;
    assign S3413 = (X[21] & Y[32]) ^ S3412;
    assign S3414 = (X[22] & Y[31]) ^ S3413;
    assign S3415 = (X[23] & Y[30]) ^ S3414;
    assign S3416 = (X[24] & Y[29]) ^ S3415;
    assign S3417 = (X[25] & Y[28]) ^ S3416;
    assign S3418 = (X[26] & Y[27]) ^ S3417;
    assign S3419 = (X[27] & Y[26]) ^ S3418;
    assign S3420 = (X[28] & Y[25]) ^ S3419;
    assign S3421 = (X[29] & Y[24]) ^ S3420;
    assign S3422 = (X[30] & Y[23]) ^ S3421;
    assign S3423 = (X[31] & Y[22]) ^ S3422;
    assign S3424 = (X[32] & Y[21]) ^ S3423;
    assign S3425 = (X[33] & Y[20]) ^ S3424;
    assign S3426 = (X[34] & Y[19]) ^ S3425;
    assign S3427 = (X[35] & Y[18]) ^ S3426;
    assign S3428 = (X[36] & Y[17]) ^ S3427;
    assign S3429 = (X[37] & Y[16]) ^ S3428;
    assign S3430 = (X[38] & Y[15]) ^ S3429;
    assign S3431 = (X[39] & Y[14]) ^ S3430;
    assign S3432 = (X[40] & Y[13]) ^ S3431;
    assign S3433 = (X[41] & Y[12]) ^ S3432;
    assign S3434 = (X[42] & Y[11]) ^ S3433;
    assign S3435 = (X[43] & Y[10]) ^ S3434;
    assign S3436 = (X[44] & Y[9]) ^ S3435;
    assign S3437 = (X[45] & Y[8]) ^ S3436;
    assign S3438 = (X[46] & Y[7]) ^ S3437;
    assign S3439 = (X[47] & Y[6]) ^ S3438;
    assign S3440 = (X[48] & Y[5]) ^ S3439;
    assign S3441 = (X[49] & Y[4]) ^ S3440;
    assign S3442 = (X[50] & Y[3]) ^ S3441;
    assign S3443 = (X[51] & Y[2]) ^ S3442;
    assign S3444 = (X[52] & Y[1]) ^ S3443;
    assign S3445 = (X[53] & Y[0]) ^ S3444;
    assign ClmulResult[53] = S3445;
    assign S3456 = X[0] & Y[54];
    assign S3457 = (X[1] & Y[53]) ^ S3456;
    assign S3458 = (X[2] & Y[52]) ^ S3457;
    assign S3459 = (X[3] & Y[51]) ^ S3458;
    assign S3460 = (X[4] & Y[50]) ^ S3459;
    assign S3461 = (X[5] & Y[49]) ^ S3460;
    assign S3462 = (X[6] & Y[48]) ^ S3461;
    assign S3463 = (X[7] & Y[47]) ^ S3462;
    assign S3464 = (X[8] & Y[46]) ^ S3463;
    assign S3465 = (X[9] & Y[45]) ^ S3464;
    assign S3466 = (X[10] & Y[44]) ^ S3465;
    assign S3467 = (X[11] & Y[43]) ^ S3466;
    assign S3468 = (X[12] & Y[42]) ^ S3467;
    assign S3469 = (X[13] & Y[41]) ^ S3468;
    assign S3470 = (X[14] & Y[40]) ^ S3469;
    assign S3471 = (X[15] & Y[39]) ^ S3470;
    assign S3472 = (X[16] & Y[38]) ^ S3471;
    assign S3473 = (X[17] & Y[37]) ^ S3472;
    assign S3474 = (X[18] & Y[36]) ^ S3473;
    assign S3475 = (X[19] & Y[35]) ^ S3474;
    assign S3476 = (X[20] & Y[34]) ^ S3475;
    assign S3477 = (X[21] & Y[33]) ^ S3476;
    assign S3478 = (X[22] & Y[32]) ^ S3477;
    assign S3479 = (X[23] & Y[31]) ^ S3478;
    assign S3480 = (X[24] & Y[30]) ^ S3479;
    assign S3481 = (X[25] & Y[29]) ^ S3480;
    assign S3482 = (X[26] & Y[28]) ^ S3481;
    assign S3483 = (X[27] & Y[27]) ^ S3482;
    assign S3484 = (X[28] & Y[26]) ^ S3483;
    assign S3485 = (X[29] & Y[25]) ^ S3484;
    assign S3486 = (X[30] & Y[24]) ^ S3485;
    assign S3487 = (X[31] & Y[23]) ^ S3486;
    assign S3488 = (X[32] & Y[22]) ^ S3487;
    assign S3489 = (X[33] & Y[21]) ^ S3488;
    assign S3490 = (X[34] & Y[20]) ^ S3489;
    assign S3491 = (X[35] & Y[19]) ^ S3490;
    assign S3492 = (X[36] & Y[18]) ^ S3491;
    assign S3493 = (X[37] & Y[17]) ^ S3492;
    assign S3494 = (X[38] & Y[16]) ^ S3493;
    assign S3495 = (X[39] & Y[15]) ^ S3494;
    assign S3496 = (X[40] & Y[14]) ^ S3495;
    assign S3497 = (X[41] & Y[13]) ^ S3496;
    assign S3498 = (X[42] & Y[12]) ^ S3497;
    assign S3499 = (X[43] & Y[11]) ^ S3498;
    assign S3500 = (X[44] & Y[10]) ^ S3499;
    assign S3501 = (X[45] & Y[9]) ^ S3500;
    assign S3502 = (X[46] & Y[8]) ^ S3501;
    assign S3503 = (X[47] & Y[7]) ^ S3502;
    assign S3504 = (X[48] & Y[6]) ^ S3503;
    assign S3505 = (X[49] & Y[5]) ^ S3504;
    assign S3506 = (X[50] & Y[4]) ^ S3505;
    assign S3507 = (X[51] & Y[3]) ^ S3506;
    assign S3508 = (X[52] & Y[2]) ^ S3507;
    assign S3509 = (X[53] & Y[1]) ^ S3508;
    assign S3510 = (X[54] & Y[0]) ^ S3509;
    assign ClmulResult[54] = S3510;
    assign S3520 = X[0] & Y[55];
    assign S3521 = (X[1] & Y[54]) ^ S3520;
    assign S3522 = (X[2] & Y[53]) ^ S3521;
    assign S3523 = (X[3] & Y[52]) ^ S3522;
    assign S3524 = (X[4] & Y[51]) ^ S3523;
    assign S3525 = (X[5] & Y[50]) ^ S3524;
    assign S3526 = (X[6] & Y[49]) ^ S3525;
    assign S3527 = (X[7] & Y[48]) ^ S3526;
    assign S3528 = (X[8] & Y[47]) ^ S3527;
    assign S3529 = (X[9] & Y[46]) ^ S3528;
    assign S3530 = (X[10] & Y[45]) ^ S3529;
    assign S3531 = (X[11] & Y[44]) ^ S3530;
    assign S3532 = (X[12] & Y[43]) ^ S3531;
    assign S3533 = (X[13] & Y[42]) ^ S3532;
    assign S3534 = (X[14] & Y[41]) ^ S3533;
    assign S3535 = (X[15] & Y[40]) ^ S3534;
    assign S3536 = (X[16] & Y[39]) ^ S3535;
    assign S3537 = (X[17] & Y[38]) ^ S3536;
    assign S3538 = (X[18] & Y[37]) ^ S3537;
    assign S3539 = (X[19] & Y[36]) ^ S3538;
    assign S3540 = (X[20] & Y[35]) ^ S3539;
    assign S3541 = (X[21] & Y[34]) ^ S3540;
    assign S3542 = (X[22] & Y[33]) ^ S3541;
    assign S3543 = (X[23] & Y[32]) ^ S3542;
    assign S3544 = (X[24] & Y[31]) ^ S3543;
    assign S3545 = (X[25] & Y[30]) ^ S3544;
    assign S3546 = (X[26] & Y[29]) ^ S3545;
    assign S3547 = (X[27] & Y[28]) ^ S3546;
    assign S3548 = (X[28] & Y[27]) ^ S3547;
    assign S3549 = (X[29] & Y[26]) ^ S3548;
    assign S3550 = (X[30] & Y[25]) ^ S3549;
    assign S3551 = (X[31] & Y[24]) ^ S3550;
    assign S3552 = (X[32] & Y[23]) ^ S3551;
    assign S3553 = (X[33] & Y[22]) ^ S3552;
    assign S3554 = (X[34] & Y[21]) ^ S3553;
    assign S3555 = (X[35] & Y[20]) ^ S3554;
    assign S3556 = (X[36] & Y[19]) ^ S3555;
    assign S3557 = (X[37] & Y[18]) ^ S3556;
    assign S3558 = (X[38] & Y[17]) ^ S3557;
    assign S3559 = (X[39] & Y[16]) ^ S3558;
    assign S3560 = (X[40] & Y[15]) ^ S3559;
    assign S3561 = (X[41] & Y[14]) ^ S3560;
    assign S3562 = (X[42] & Y[13]) ^ S3561;
    assign S3563 = (X[43] & Y[12]) ^ S3562;
    assign S3564 = (X[44] & Y[11]) ^ S3563;
    assign S3565 = (X[45] & Y[10]) ^ S3564;
    assign S3566 = (X[46] & Y[9]) ^ S3565;
    assign S3567 = (X[47] & Y[8]) ^ S3566;
    assign S3568 = (X[48] & Y[7]) ^ S3567;
    assign S3569 = (X[49] & Y[6]) ^ S3568;
    assign S3570 = (X[50] & Y[5]) ^ S3569;
    assign S3571 = (X[51] & Y[4]) ^ S3570;
    assign S3572 = (X[52] & Y[3]) ^ S3571;
    assign S3573 = (X[53] & Y[2]) ^ S3572;
    assign S3574 = (X[54] & Y[1]) ^ S3573;
    assign S3575 = (X[55] & Y[0]) ^ S3574;
    assign ClmulResult[55] = S3575;
    assign S3584 = X[0] & Y[56];
    assign S3585 = (X[1] & Y[55]) ^ S3584;
    assign S3586 = (X[2] & Y[54]) ^ S3585;
    assign S3587 = (X[3] & Y[53]) ^ S3586;
    assign S3588 = (X[4] & Y[52]) ^ S3587;
    assign S3589 = (X[5] & Y[51]) ^ S3588;
    assign S3590 = (X[6] & Y[50]) ^ S3589;
    assign S3591 = (X[7] & Y[49]) ^ S3590;
    assign S3592 = (X[8] & Y[48]) ^ S3591;
    assign S3593 = (X[9] & Y[47]) ^ S3592;
    assign S3594 = (X[10] & Y[46]) ^ S3593;
    assign S3595 = (X[11] & Y[45]) ^ S3594;
    assign S3596 = (X[12] & Y[44]) ^ S3595;
    assign S3597 = (X[13] & Y[43]) ^ S3596;
    assign S3598 = (X[14] & Y[42]) ^ S3597;
    assign S3599 = (X[15] & Y[41]) ^ S3598;
    assign S3600 = (X[16] & Y[40]) ^ S3599;
    assign S3601 = (X[17] & Y[39]) ^ S3600;
    assign S3602 = (X[18] & Y[38]) ^ S3601;
    assign S3603 = (X[19] & Y[37]) ^ S3602;
    assign S3604 = (X[20] & Y[36]) ^ S3603;
    assign S3605 = (X[21] & Y[35]) ^ S3604;
    assign S3606 = (X[22] & Y[34]) ^ S3605;
    assign S3607 = (X[23] & Y[33]) ^ S3606;
    assign S3608 = (X[24] & Y[32]) ^ S3607;
    assign S3609 = (X[25] & Y[31]) ^ S3608;
    assign S3610 = (X[26] & Y[30]) ^ S3609;
    assign S3611 = (X[27] & Y[29]) ^ S3610;
    assign S3612 = (X[28] & Y[28]) ^ S3611;
    assign S3613 = (X[29] & Y[27]) ^ S3612;
    assign S3614 = (X[30] & Y[26]) ^ S3613;
    assign S3615 = (X[31] & Y[25]) ^ S3614;
    assign S3616 = (X[32] & Y[24]) ^ S3615;
    assign S3617 = (X[33] & Y[23]) ^ S3616;
    assign S3618 = (X[34] & Y[22]) ^ S3617;
    assign S3619 = (X[35] & Y[21]) ^ S3618;
    assign S3620 = (X[36] & Y[20]) ^ S3619;
    assign S3621 = (X[37] & Y[19]) ^ S3620;
    assign S3622 = (X[38] & Y[18]) ^ S3621;
    assign S3623 = (X[39] & Y[17]) ^ S3622;
    assign S3624 = (X[40] & Y[16]) ^ S3623;
    assign S3625 = (X[41] & Y[15]) ^ S3624;
    assign S3626 = (X[42] & Y[14]) ^ S3625;
    assign S3627 = (X[43] & Y[13]) ^ S3626;
    assign S3628 = (X[44] & Y[12]) ^ S3627;
    assign S3629 = (X[45] & Y[11]) ^ S3628;
    assign S3630 = (X[46] & Y[10]) ^ S3629;
    assign S3631 = (X[47] & Y[9]) ^ S3630;
    assign S3632 = (X[48] & Y[8]) ^ S3631;
    assign S3633 = (X[49] & Y[7]) ^ S3632;
    assign S3634 = (X[50] & Y[6]) ^ S3633;
    assign S3635 = (X[51] & Y[5]) ^ S3634;
    assign S3636 = (X[52] & Y[4]) ^ S3635;
    assign S3637 = (X[53] & Y[3]) ^ S3636;
    assign S3638 = (X[54] & Y[2]) ^ S3637;
    assign S3639 = (X[55] & Y[1]) ^ S3638;
    assign S3640 = (X[56] & Y[0]) ^ S3639;
    assign ClmulResult[56] = S3640;
    assign S3648 = X[0] & Y[57];
    assign S3649 = (X[1] & Y[56]) ^ S3648;
    assign S3650 = (X[2] & Y[55]) ^ S3649;
    assign S3651 = (X[3] & Y[54]) ^ S3650;
    assign S3652 = (X[4] & Y[53]) ^ S3651;
    assign S3653 = (X[5] & Y[52]) ^ S3652;
    assign S3654 = (X[6] & Y[51]) ^ S3653;
    assign S3655 = (X[7] & Y[50]) ^ S3654;
    assign S3656 = (X[8] & Y[49]) ^ S3655;
    assign S3657 = (X[9] & Y[48]) ^ S3656;
    assign S3658 = (X[10] & Y[47]) ^ S3657;
    assign S3659 = (X[11] & Y[46]) ^ S3658;
    assign S3660 = (X[12] & Y[45]) ^ S3659;
    assign S3661 = (X[13] & Y[44]) ^ S3660;
    assign S3662 = (X[14] & Y[43]) ^ S3661;
    assign S3663 = (X[15] & Y[42]) ^ S3662;
    assign S3664 = (X[16] & Y[41]) ^ S3663;
    assign S3665 = (X[17] & Y[40]) ^ S3664;
    assign S3666 = (X[18] & Y[39]) ^ S3665;
    assign S3667 = (X[19] & Y[38]) ^ S3666;
    assign S3668 = (X[20] & Y[37]) ^ S3667;
    assign S3669 = (X[21] & Y[36]) ^ S3668;
    assign S3670 = (X[22] & Y[35]) ^ S3669;
    assign S3671 = (X[23] & Y[34]) ^ S3670;
    assign S3672 = (X[24] & Y[33]) ^ S3671;
    assign S3673 = (X[25] & Y[32]) ^ S3672;
    assign S3674 = (X[26] & Y[31]) ^ S3673;
    assign S3675 = (X[27] & Y[30]) ^ S3674;
    assign S3676 = (X[28] & Y[29]) ^ S3675;
    assign S3677 = (X[29] & Y[28]) ^ S3676;
    assign S3678 = (X[30] & Y[27]) ^ S3677;
    assign S3679 = (X[31] & Y[26]) ^ S3678;
    assign S3680 = (X[32] & Y[25]) ^ S3679;
    assign S3681 = (X[33] & Y[24]) ^ S3680;
    assign S3682 = (X[34] & Y[23]) ^ S3681;
    assign S3683 = (X[35] & Y[22]) ^ S3682;
    assign S3684 = (X[36] & Y[21]) ^ S3683;
    assign S3685 = (X[37] & Y[20]) ^ S3684;
    assign S3686 = (X[38] & Y[19]) ^ S3685;
    assign S3687 = (X[39] & Y[18]) ^ S3686;
    assign S3688 = (X[40] & Y[17]) ^ S3687;
    assign S3689 = (X[41] & Y[16]) ^ S3688;
    assign S3690 = (X[42] & Y[15]) ^ S3689;
    assign S3691 = (X[43] & Y[14]) ^ S3690;
    assign S3692 = (X[44] & Y[13]) ^ S3691;
    assign S3693 = (X[45] & Y[12]) ^ S3692;
    assign S3694 = (X[46] & Y[11]) ^ S3693;
    assign S3695 = (X[47] & Y[10]) ^ S3694;
    assign S3696 = (X[48] & Y[9]) ^ S3695;
    assign S3697 = (X[49] & Y[8]) ^ S3696;
    assign S3698 = (X[50] & Y[7]) ^ S3697;
    assign S3699 = (X[51] & Y[6]) ^ S3698;
    assign S3700 = (X[52] & Y[5]) ^ S3699;
    assign S3701 = (X[53] & Y[4]) ^ S3700;
    assign S3702 = (X[54] & Y[3]) ^ S3701;
    assign S3703 = (X[55] & Y[2]) ^ S3702;
    assign S3704 = (X[56] & Y[1]) ^ S3703;
    assign S3705 = (X[57] & Y[0]) ^ S3704;
    assign ClmulResult[57] = S3705;
    assign S3712 = X[0] & Y[58];
    assign S3713 = (X[1] & Y[57]) ^ S3712;
    assign S3714 = (X[2] & Y[56]) ^ S3713;
    assign S3715 = (X[3] & Y[55]) ^ S3714;
    assign S3716 = (X[4] & Y[54]) ^ S3715;
    assign S3717 = (X[5] & Y[53]) ^ S3716;
    assign S3718 = (X[6] & Y[52]) ^ S3717;
    assign S3719 = (X[7] & Y[51]) ^ S3718;
    assign S3720 = (X[8] & Y[50]) ^ S3719;
    assign S3721 = (X[9] & Y[49]) ^ S3720;
    assign S3722 = (X[10] & Y[48]) ^ S3721;
    assign S3723 = (X[11] & Y[47]) ^ S3722;
    assign S3724 = (X[12] & Y[46]) ^ S3723;
    assign S3725 = (X[13] & Y[45]) ^ S3724;
    assign S3726 = (X[14] & Y[44]) ^ S3725;
    assign S3727 = (X[15] & Y[43]) ^ S3726;
    assign S3728 = (X[16] & Y[42]) ^ S3727;
    assign S3729 = (X[17] & Y[41]) ^ S3728;
    assign S3730 = (X[18] & Y[40]) ^ S3729;
    assign S3731 = (X[19] & Y[39]) ^ S3730;
    assign S3732 = (X[20] & Y[38]) ^ S3731;
    assign S3733 = (X[21] & Y[37]) ^ S3732;
    assign S3734 = (X[22] & Y[36]) ^ S3733;
    assign S3735 = (X[23] & Y[35]) ^ S3734;
    assign S3736 = (X[24] & Y[34]) ^ S3735;
    assign S3737 = (X[25] & Y[33]) ^ S3736;
    assign S3738 = (X[26] & Y[32]) ^ S3737;
    assign S3739 = (X[27] & Y[31]) ^ S3738;
    assign S3740 = (X[28] & Y[30]) ^ S3739;
    assign S3741 = (X[29] & Y[29]) ^ S3740;
    assign S3742 = (X[30] & Y[28]) ^ S3741;
    assign S3743 = (X[31] & Y[27]) ^ S3742;
    assign S3744 = (X[32] & Y[26]) ^ S3743;
    assign S3745 = (X[33] & Y[25]) ^ S3744;
    assign S3746 = (X[34] & Y[24]) ^ S3745;
    assign S3747 = (X[35] & Y[23]) ^ S3746;
    assign S3748 = (X[36] & Y[22]) ^ S3747;
    assign S3749 = (X[37] & Y[21]) ^ S3748;
    assign S3750 = (X[38] & Y[20]) ^ S3749;
    assign S3751 = (X[39] & Y[19]) ^ S3750;
    assign S3752 = (X[40] & Y[18]) ^ S3751;
    assign S3753 = (X[41] & Y[17]) ^ S3752;
    assign S3754 = (X[42] & Y[16]) ^ S3753;
    assign S3755 = (X[43] & Y[15]) ^ S3754;
    assign S3756 = (X[44] & Y[14]) ^ S3755;
    assign S3757 = (X[45] & Y[13]) ^ S3756;
    assign S3758 = (X[46] & Y[12]) ^ S3757;
    assign S3759 = (X[47] & Y[11]) ^ S3758;
    assign S3760 = (X[48] & Y[10]) ^ S3759;
    assign S3761 = (X[49] & Y[9]) ^ S3760;
    assign S3762 = (X[50] & Y[8]) ^ S3761;
    assign S3763 = (X[51] & Y[7]) ^ S3762;
    assign S3764 = (X[52] & Y[6]) ^ S3763;
    assign S3765 = (X[53] & Y[5]) ^ S3764;
    assign S3766 = (X[54] & Y[4]) ^ S3765;
    assign S3767 = (X[55] & Y[3]) ^ S3766;
    assign S3768 = (X[56] & Y[2]) ^ S3767;
    assign S3769 = (X[57] & Y[1]) ^ S3768;
    assign S3770 = (X[58] & Y[0]) ^ S3769;
    assign ClmulResult[58] = S3770;
    assign S3776 = X[0] & Y[59];
    assign S3777 = (X[1] & Y[58]) ^ S3776;
    assign S3778 = (X[2] & Y[57]) ^ S3777;
    assign S3779 = (X[3] & Y[56]) ^ S3778;
    assign S3780 = (X[4] & Y[55]) ^ S3779;
    assign S3781 = (X[5] & Y[54]) ^ S3780;
    assign S3782 = (X[6] & Y[53]) ^ S3781;
    assign S3783 = (X[7] & Y[52]) ^ S3782;
    assign S3784 = (X[8] & Y[51]) ^ S3783;
    assign S3785 = (X[9] & Y[50]) ^ S3784;
    assign S3786 = (X[10] & Y[49]) ^ S3785;
    assign S3787 = (X[11] & Y[48]) ^ S3786;
    assign S3788 = (X[12] & Y[47]) ^ S3787;
    assign S3789 = (X[13] & Y[46]) ^ S3788;
    assign S3790 = (X[14] & Y[45]) ^ S3789;
    assign S3791 = (X[15] & Y[44]) ^ S3790;
    assign S3792 = (X[16] & Y[43]) ^ S3791;
    assign S3793 = (X[17] & Y[42]) ^ S3792;
    assign S3794 = (X[18] & Y[41]) ^ S3793;
    assign S3795 = (X[19] & Y[40]) ^ S3794;
    assign S3796 = (X[20] & Y[39]) ^ S3795;
    assign S3797 = (X[21] & Y[38]) ^ S3796;
    assign S3798 = (X[22] & Y[37]) ^ S3797;
    assign S3799 = (X[23] & Y[36]) ^ S3798;
    assign S3800 = (X[24] & Y[35]) ^ S3799;
    assign S3801 = (X[25] & Y[34]) ^ S3800;
    assign S3802 = (X[26] & Y[33]) ^ S3801;
    assign S3803 = (X[27] & Y[32]) ^ S3802;
    assign S3804 = (X[28] & Y[31]) ^ S3803;
    assign S3805 = (X[29] & Y[30]) ^ S3804;
    assign S3806 = (X[30] & Y[29]) ^ S3805;
    assign S3807 = (X[31] & Y[28]) ^ S3806;
    assign S3808 = (X[32] & Y[27]) ^ S3807;
    assign S3809 = (X[33] & Y[26]) ^ S3808;
    assign S3810 = (X[34] & Y[25]) ^ S3809;
    assign S3811 = (X[35] & Y[24]) ^ S3810;
    assign S3812 = (X[36] & Y[23]) ^ S3811;
    assign S3813 = (X[37] & Y[22]) ^ S3812;
    assign S3814 = (X[38] & Y[21]) ^ S3813;
    assign S3815 = (X[39] & Y[20]) ^ S3814;
    assign S3816 = (X[40] & Y[19]) ^ S3815;
    assign S3817 = (X[41] & Y[18]) ^ S3816;
    assign S3818 = (X[42] & Y[17]) ^ S3817;
    assign S3819 = (X[43] & Y[16]) ^ S3818;
    assign S3820 = (X[44] & Y[15]) ^ S3819;
    assign S3821 = (X[45] & Y[14]) ^ S3820;
    assign S3822 = (X[46] & Y[13]) ^ S3821;
    assign S3823 = (X[47] & Y[12]) ^ S3822;
    assign S3824 = (X[48] & Y[11]) ^ S3823;
    assign S3825 = (X[49] & Y[10]) ^ S3824;
    assign S3826 = (X[50] & Y[9]) ^ S3825;
    assign S3827 = (X[51] & Y[8]) ^ S3826;
    assign S3828 = (X[52] & Y[7]) ^ S3827;
    assign S3829 = (X[53] & Y[6]) ^ S3828;
    assign S3830 = (X[54] & Y[5]) ^ S3829;
    assign S3831 = (X[55] & Y[4]) ^ S3830;
    assign S3832 = (X[56] & Y[3]) ^ S3831;
    assign S3833 = (X[57] & Y[2]) ^ S3832;
    assign S3834 = (X[58] & Y[1]) ^ S3833;
    assign S3835 = (X[59] & Y[0]) ^ S3834;
    assign ClmulResult[59] = S3835;
    assign S3840 = X[0] & Y[60];
    assign S3841 = (X[1] & Y[59]) ^ S3840;
    assign S3842 = (X[2] & Y[58]) ^ S3841;
    assign S3843 = (X[3] & Y[57]) ^ S3842;
    assign S3844 = (X[4] & Y[56]) ^ S3843;
    assign S3845 = (X[5] & Y[55]) ^ S3844;
    assign S3846 = (X[6] & Y[54]) ^ S3845;
    assign S3847 = (X[7] & Y[53]) ^ S3846;
    assign S3848 = (X[8] & Y[52]) ^ S3847;
    assign S3849 = (X[9] & Y[51]) ^ S3848;
    assign S3850 = (X[10] & Y[50]) ^ S3849;
    assign S3851 = (X[11] & Y[49]) ^ S3850;
    assign S3852 = (X[12] & Y[48]) ^ S3851;
    assign S3853 = (X[13] & Y[47]) ^ S3852;
    assign S3854 = (X[14] & Y[46]) ^ S3853;
    assign S3855 = (X[15] & Y[45]) ^ S3854;
    assign S3856 = (X[16] & Y[44]) ^ S3855;
    assign S3857 = (X[17] & Y[43]) ^ S3856;
    assign S3858 = (X[18] & Y[42]) ^ S3857;
    assign S3859 = (X[19] & Y[41]) ^ S3858;
    assign S3860 = (X[20] & Y[40]) ^ S3859;
    assign S3861 = (X[21] & Y[39]) ^ S3860;
    assign S3862 = (X[22] & Y[38]) ^ S3861;
    assign S3863 = (X[23] & Y[37]) ^ S3862;
    assign S3864 = (X[24] & Y[36]) ^ S3863;
    assign S3865 = (X[25] & Y[35]) ^ S3864;
    assign S3866 = (X[26] & Y[34]) ^ S3865;
    assign S3867 = (X[27] & Y[33]) ^ S3866;
    assign S3868 = (X[28] & Y[32]) ^ S3867;
    assign S3869 = (X[29] & Y[31]) ^ S3868;
    assign S3870 = (X[30] & Y[30]) ^ S3869;
    assign S3871 = (X[31] & Y[29]) ^ S3870;
    assign S3872 = (X[32] & Y[28]) ^ S3871;
    assign S3873 = (X[33] & Y[27]) ^ S3872;
    assign S3874 = (X[34] & Y[26]) ^ S3873;
    assign S3875 = (X[35] & Y[25]) ^ S3874;
    assign S3876 = (X[36] & Y[24]) ^ S3875;
    assign S3877 = (X[37] & Y[23]) ^ S3876;
    assign S3878 = (X[38] & Y[22]) ^ S3877;
    assign S3879 = (X[39] & Y[21]) ^ S3878;
    assign S3880 = (X[40] & Y[20]) ^ S3879;
    assign S3881 = (X[41] & Y[19]) ^ S3880;
    assign S3882 = (X[42] & Y[18]) ^ S3881;
    assign S3883 = (X[43] & Y[17]) ^ S3882;
    assign S3884 = (X[44] & Y[16]) ^ S3883;
    assign S3885 = (X[45] & Y[15]) ^ S3884;
    assign S3886 = (X[46] & Y[14]) ^ S3885;
    assign S3887 = (X[47] & Y[13]) ^ S3886;
    assign S3888 = (X[48] & Y[12]) ^ S3887;
    assign S3889 = (X[49] & Y[11]) ^ S3888;
    assign S3890 = (X[50] & Y[10]) ^ S3889;
    assign S3891 = (X[51] & Y[9]) ^ S3890;
    assign S3892 = (X[52] & Y[8]) ^ S3891;
    assign S3893 = (X[53] & Y[7]) ^ S3892;
    assign S3894 = (X[54] & Y[6]) ^ S3893;
    assign S3895 = (X[55] & Y[5]) ^ S3894;
    assign S3896 = (X[56] & Y[4]) ^ S3895;
    assign S3897 = (X[57] & Y[3]) ^ S3896;
    assign S3898 = (X[58] & Y[2]) ^ S3897;
    assign S3899 = (X[59] & Y[1]) ^ S3898;
    assign S3900 = (X[60] & Y[0]) ^ S3899;
    assign ClmulResult[60] = S3900;
    assign S3904 = X[0] & Y[61];
    assign S3905 = (X[1] & Y[60]) ^ S3904;
    assign S3906 = (X[2] & Y[59]) ^ S3905;
    assign S3907 = (X[3] & Y[58]) ^ S3906;
    assign S3908 = (X[4] & Y[57]) ^ S3907;
    assign S3909 = (X[5] & Y[56]) ^ S3908;
    assign S3910 = (X[6] & Y[55]) ^ S3909;
    assign S3911 = (X[7] & Y[54]) ^ S3910;
    assign S3912 = (X[8] & Y[53]) ^ S3911;
    assign S3913 = (X[9] & Y[52]) ^ S3912;
    assign S3914 = (X[10] & Y[51]) ^ S3913;
    assign S3915 = (X[11] & Y[50]) ^ S3914;
    assign S3916 = (X[12] & Y[49]) ^ S3915;
    assign S3917 = (X[13] & Y[48]) ^ S3916;
    assign S3918 = (X[14] & Y[47]) ^ S3917;
    assign S3919 = (X[15] & Y[46]) ^ S3918;
    assign S3920 = (X[16] & Y[45]) ^ S3919;
    assign S3921 = (X[17] & Y[44]) ^ S3920;
    assign S3922 = (X[18] & Y[43]) ^ S3921;
    assign S3923 = (X[19] & Y[42]) ^ S3922;
    assign S3924 = (X[20] & Y[41]) ^ S3923;
    assign S3925 = (X[21] & Y[40]) ^ S3924;
    assign S3926 = (X[22] & Y[39]) ^ S3925;
    assign S3927 = (X[23] & Y[38]) ^ S3926;
    assign S3928 = (X[24] & Y[37]) ^ S3927;
    assign S3929 = (X[25] & Y[36]) ^ S3928;
    assign S3930 = (X[26] & Y[35]) ^ S3929;
    assign S3931 = (X[27] & Y[34]) ^ S3930;
    assign S3932 = (X[28] & Y[33]) ^ S3931;
    assign S3933 = (X[29] & Y[32]) ^ S3932;
    assign S3934 = (X[30] & Y[31]) ^ S3933;
    assign S3935 = (X[31] & Y[30]) ^ S3934;
    assign S3936 = (X[32] & Y[29]) ^ S3935;
    assign S3937 = (X[33] & Y[28]) ^ S3936;
    assign S3938 = (X[34] & Y[27]) ^ S3937;
    assign S3939 = (X[35] & Y[26]) ^ S3938;
    assign S3940 = (X[36] & Y[25]) ^ S3939;
    assign S3941 = (X[37] & Y[24]) ^ S3940;
    assign S3942 = (X[38] & Y[23]) ^ S3941;
    assign S3943 = (X[39] & Y[22]) ^ S3942;
    assign S3944 = (X[40] & Y[21]) ^ S3943;
    assign S3945 = (X[41] & Y[20]) ^ S3944;
    assign S3946 = (X[42] & Y[19]) ^ S3945;
    assign S3947 = (X[43] & Y[18]) ^ S3946;
    assign S3948 = (X[44] & Y[17]) ^ S3947;
    assign S3949 = (X[45] & Y[16]) ^ S3948;
    assign S3950 = (X[46] & Y[15]) ^ S3949;
    assign S3951 = (X[47] & Y[14]) ^ S3950;
    assign S3952 = (X[48] & Y[13]) ^ S3951;
    assign S3953 = (X[49] & Y[12]) ^ S3952;
    assign S3954 = (X[50] & Y[11]) ^ S3953;
    assign S3955 = (X[51] & Y[10]) ^ S3954;
    assign S3956 = (X[52] & Y[9]) ^ S3955;
    assign S3957 = (X[53] & Y[8]) ^ S3956;
    assign S3958 = (X[54] & Y[7]) ^ S3957;
    assign S3959 = (X[55] & Y[6]) ^ S3958;
    assign S3960 = (X[56] & Y[5]) ^ S3959;
    assign S3961 = (X[57] & Y[4]) ^ S3960;
    assign S3962 = (X[58] & Y[3]) ^ S3961;
    assign S3963 = (X[59] & Y[2]) ^ S3962;
    assign S3964 = (X[60] & Y[1]) ^ S3963;
    assign S3965 = (X[61] & Y[0]) ^ S3964;
    assign ClmulResult[61] = S3965;
    assign S3968 = X[0] & Y[62];
    assign S3969 = (X[1] & Y[61]) ^ S3968;
    assign S3970 = (X[2] & Y[60]) ^ S3969;
    assign S3971 = (X[3] & Y[59]) ^ S3970;
    assign S3972 = (X[4] & Y[58]) ^ S3971;
    assign S3973 = (X[5] & Y[57]) ^ S3972;
    assign S3974 = (X[6] & Y[56]) ^ S3973;
    assign S3975 = (X[7] & Y[55]) ^ S3974;
    assign S3976 = (X[8] & Y[54]) ^ S3975;
    assign S3977 = (X[9] & Y[53]) ^ S3976;
    assign S3978 = (X[10] & Y[52]) ^ S3977;
    assign S3979 = (X[11] & Y[51]) ^ S3978;
    assign S3980 = (X[12] & Y[50]) ^ S3979;
    assign S3981 = (X[13] & Y[49]) ^ S3980;
    assign S3982 = (X[14] & Y[48]) ^ S3981;
    assign S3983 = (X[15] & Y[47]) ^ S3982;
    assign S3984 = (X[16] & Y[46]) ^ S3983;
    assign S3985 = (X[17] & Y[45]) ^ S3984;
    assign S3986 = (X[18] & Y[44]) ^ S3985;
    assign S3987 = (X[19] & Y[43]) ^ S3986;
    assign S3988 = (X[20] & Y[42]) ^ S3987;
    assign S3989 = (X[21] & Y[41]) ^ S3988;
    assign S3990 = (X[22] & Y[40]) ^ S3989;
    assign S3991 = (X[23] & Y[39]) ^ S3990;
    assign S3992 = (X[24] & Y[38]) ^ S3991;
    assign S3993 = (X[25] & Y[37]) ^ S3992;
    assign S3994 = (X[26] & Y[36]) ^ S3993;
    assign S3995 = (X[27] & Y[35]) ^ S3994;
    assign S3996 = (X[28] & Y[34]) ^ S3995;
    assign S3997 = (X[29] & Y[33]) ^ S3996;
    assign S3998 = (X[30] & Y[32]) ^ S3997;
    assign S3999 = (X[31] & Y[31]) ^ S3998;
    assign S4000 = (X[32] & Y[30]) ^ S3999;
    assign S4001 = (X[33] & Y[29]) ^ S4000;
    assign S4002 = (X[34] & Y[28]) ^ S4001;
    assign S4003 = (X[35] & Y[27]) ^ S4002;
    assign S4004 = (X[36] & Y[26]) ^ S4003;
    assign S4005 = (X[37] & Y[25]) ^ S4004;
    assign S4006 = (X[38] & Y[24]) ^ S4005;
    assign S4007 = (X[39] & Y[23]) ^ S4006;
    assign S4008 = (X[40] & Y[22]) ^ S4007;
    assign S4009 = (X[41] & Y[21]) ^ S4008;
    assign S4010 = (X[42] & Y[20]) ^ S4009;
    assign S4011 = (X[43] & Y[19]) ^ S4010;
    assign S4012 = (X[44] & Y[18]) ^ S4011;
    assign S4013 = (X[45] & Y[17]) ^ S4012;
    assign S4014 = (X[46] & Y[16]) ^ S4013;
    assign S4015 = (X[47] & Y[15]) ^ S4014;
    assign S4016 = (X[48] & Y[14]) ^ S4015;
    assign S4017 = (X[49] & Y[13]) ^ S4016;
    assign S4018 = (X[50] & Y[12]) ^ S4017;
    assign S4019 = (X[51] & Y[11]) ^ S4018;
    assign S4020 = (X[52] & Y[10]) ^ S4019;
    assign S4021 = (X[53] & Y[9]) ^ S4020;
    assign S4022 = (X[54] & Y[8]) ^ S4021;
    assign S4023 = (X[55] & Y[7]) ^ S4022;
    assign S4024 = (X[56] & Y[6]) ^ S4023;
    assign S4025 = (X[57] & Y[5]) ^ S4024;
    assign S4026 = (X[58] & Y[4]) ^ S4025;
    assign S4027 = (X[59] & Y[3]) ^ S4026;
    assign S4028 = (X[60] & Y[2]) ^ S4027;
    assign S4029 = (X[61] & Y[1]) ^ S4028;
    assign S4030 = (X[62] & Y[0]) ^ S4029;
    assign ClmulResult[62] = S4030;
    assign S4032 = X[0] & Y[63];
    assign S4033 = (X[1] & Y[62]) ^ S4032;
    assign S4034 = (X[2] & Y[61]) ^ S4033;
    assign S4035 = (X[3] & Y[60]) ^ S4034;
    assign S4036 = (X[4] & Y[59]) ^ S4035;
    assign S4037 = (X[5] & Y[58]) ^ S4036;
    assign S4038 = (X[6] & Y[57]) ^ S4037;
    assign S4039 = (X[7] & Y[56]) ^ S4038;
    assign S4040 = (X[8] & Y[55]) ^ S4039;
    assign S4041 = (X[9] & Y[54]) ^ S4040;
    assign S4042 = (X[10] & Y[53]) ^ S4041;
    assign S4043 = (X[11] & Y[52]) ^ S4042;
    assign S4044 = (X[12] & Y[51]) ^ S4043;
    assign S4045 = (X[13] & Y[50]) ^ S4044;
    assign S4046 = (X[14] & Y[49]) ^ S4045;
    assign S4047 = (X[15] & Y[48]) ^ S4046;
    assign S4048 = (X[16] & Y[47]) ^ S4047;
    assign S4049 = (X[17] & Y[46]) ^ S4048;
    assign S4050 = (X[18] & Y[45]) ^ S4049;
    assign S4051 = (X[19] & Y[44]) ^ S4050;
    assign S4052 = (X[20] & Y[43]) ^ S4051;
    assign S4053 = (X[21] & Y[42]) ^ S4052;
    assign S4054 = (X[22] & Y[41]) ^ S4053;
    assign S4055 = (X[23] & Y[40]) ^ S4054;
    assign S4056 = (X[24] & Y[39]) ^ S4055;
    assign S4057 = (X[25] & Y[38]) ^ S4056;
    assign S4058 = (X[26] & Y[37]) ^ S4057;
    assign S4059 = (X[27] & Y[36]) ^ S4058;
    assign S4060 = (X[28] & Y[35]) ^ S4059;
    assign S4061 = (X[29] & Y[34]) ^ S4060;
    assign S4062 = (X[30] & Y[33]) ^ S4061;
    assign S4063 = (X[31] & Y[32]) ^ S4062;
    assign S4064 = (X[32] & Y[31]) ^ S4063;
    assign S4065 = (X[33] & Y[30]) ^ S4064;
    assign S4066 = (X[34] & Y[29]) ^ S4065;
    assign S4067 = (X[35] & Y[28]) ^ S4066;
    assign S4068 = (X[36] & Y[27]) ^ S4067;
    assign S4069 = (X[37] & Y[26]) ^ S4068;
    assign S4070 = (X[38] & Y[25]) ^ S4069;
    assign S4071 = (X[39] & Y[24]) ^ S4070;
    assign S4072 = (X[40] & Y[23]) ^ S4071;
    assign S4073 = (X[41] & Y[22]) ^ S4072;
    assign S4074 = (X[42] & Y[21]) ^ S4073;
    assign S4075 = (X[43] & Y[20]) ^ S4074;
    assign S4076 = (X[44] & Y[19]) ^ S4075;
    assign S4077 = (X[45] & Y[18]) ^ S4076;
    assign S4078 = (X[46] & Y[17]) ^ S4077;
    assign S4079 = (X[47] & Y[16]) ^ S4078;
    assign S4080 = (X[48] & Y[15]) ^ S4079;
    assign S4081 = (X[49] & Y[14]) ^ S4080;
    assign S4082 = (X[50] & Y[13]) ^ S4081;
    assign S4083 = (X[51] & Y[12]) ^ S4082;
    assign S4084 = (X[52] & Y[11]) ^ S4083;
    assign S4085 = (X[53] & Y[10]) ^ S4084;
    assign S4086 = (X[54] & Y[9]) ^ S4085;
    assign S4087 = (X[55] & Y[8]) ^ S4086;
    assign S4088 = (X[56] & Y[7]) ^ S4087;
    assign S4089 = (X[57] & Y[6]) ^ S4088;
    assign S4090 = (X[58] & Y[5]) ^ S4089;
    assign S4091 = (X[59] & Y[4]) ^ S4090;
    assign S4092 = (X[60] & Y[3]) ^ S4091;
    assign S4093 = (X[61] & Y[2]) ^ S4092;
    assign S4094 = (X[62] & Y[1]) ^ S4093;
    assign S4095 = (X[63] & Y[0]) ^ S4094;
    assign ClmulResult[63] = S4095;

  end
  else begin
    assign S0 = X[0] & Y[0];
    assign ClmulResult[0] = S0;
    assign S32 = X[0] & Y[1];
    assign S33 = (X[1] & Y[0]) ^ S32;
    assign ClmulResult[1] = S33;
    assign S64 = X[0] & Y[2];
    assign S65 = (X[1] & Y[1]) ^ S64;
    assign S66 = (X[2] & Y[0]) ^ S65;
    assign ClmulResult[2] = S66;
    assign S96 = X[0] & Y[3];
    assign S97 = (X[1] & Y[2]) ^ S96;
    assign S98 = (X[2] & Y[1]) ^ S97;
    assign S99 = (X[3] & Y[0]) ^ S98;
    assign ClmulResult[3] = S99;
    assign S128 = X[0] & Y[4];
    assign S129 = (X[1] & Y[3]) ^ S128;
    assign S130 = (X[2] & Y[2]) ^ S129;
    assign S131 = (X[3] & Y[1]) ^ S130;
    assign S132 = (X[4] & Y[0]) ^ S131;
    assign ClmulResult[4] = S132;
    assign S160 = X[0] & Y[5];
    assign S161 = (X[1] & Y[4]) ^ S160;
    assign S162 = (X[2] & Y[3]) ^ S161;
    assign S163 = (X[3] & Y[2]) ^ S162;
    assign S164 = (X[4] & Y[1]) ^ S163;
    assign S165 = (X[5] & Y[0]) ^ S164;
    assign ClmulResult[5] = S165;
    assign S192 = X[0] & Y[6];
    assign S193 = (X[1] & Y[5]) ^ S192;
    assign S194 = (X[2] & Y[4]) ^ S193;
    assign S195 = (X[3] & Y[3]) ^ S194;
    assign S196 = (X[4] & Y[2]) ^ S195;
    assign S197 = (X[5] & Y[1]) ^ S196;
    assign S198 = (X[6] & Y[0]) ^ S197;
    assign ClmulResult[6] = S198;
    assign S224 = X[0] & Y[7];
    assign S225 = (X[1] & Y[6]) ^ S224;
    assign S226 = (X[2] & Y[5]) ^ S225;
    assign S227 = (X[3] & Y[4]) ^ S226;
    assign S228 = (X[4] & Y[3]) ^ S227;
    assign S229 = (X[5] & Y[2]) ^ S228;
    assign S230 = (X[6] & Y[1]) ^ S229;
    assign S231 = (X[7] & Y[0]) ^ S230;
    assign ClmulResult[7] = S231;
    assign S256 = X[0] & Y[8];
    assign S257 = (X[1] & Y[7]) ^ S256;
    assign S258 = (X[2] & Y[6]) ^ S257;
    assign S259 = (X[3] & Y[5]) ^ S258;
    assign S260 = (X[4] & Y[4]) ^ S259;
    assign S261 = (X[5] & Y[3]) ^ S260;
    assign S262 = (X[6] & Y[2]) ^ S261;
    assign S263 = (X[7] & Y[1]) ^ S262;
    assign S264 = (X[8] & Y[0]) ^ S263;
    assign ClmulResult[8] = S264;
    assign S288 = X[0] & Y[9];
    assign S289 = (X[1] & Y[8]) ^ S288;
    assign S290 = (X[2] & Y[7]) ^ S289;
    assign S291 = (X[3] & Y[6]) ^ S290;
    assign S292 = (X[4] & Y[5]) ^ S291;
    assign S293 = (X[5] & Y[4]) ^ S292;
    assign S294 = (X[6] & Y[3]) ^ S293;
    assign S295 = (X[7] & Y[2]) ^ S294;
    assign S296 = (X[8] & Y[1]) ^ S295;
    assign S297 = (X[9] & Y[0]) ^ S296;
    assign ClmulResult[9] = S297;
    assign S320 = X[0] & Y[10];
    assign S321 = (X[1] & Y[9]) ^ S320;
    assign S322 = (X[2] & Y[8]) ^ S321;
    assign S323 = (X[3] & Y[7]) ^ S322;
    assign S324 = (X[4] & Y[6]) ^ S323;
    assign S325 = (X[5] & Y[5]) ^ S324;
    assign S326 = (X[6] & Y[4]) ^ S325;
    assign S327 = (X[7] & Y[3]) ^ S326;
    assign S328 = (X[8] & Y[2]) ^ S327;
    assign S329 = (X[9] & Y[1]) ^ S328;
    assign S330 = (X[10] & Y[0]) ^ S329;
    assign ClmulResult[10] = S330;
    assign S352 = X[0] & Y[11];
    assign S353 = (X[1] & Y[10]) ^ S352;
    assign S354 = (X[2] & Y[9]) ^ S353;
    assign S355 = (X[3] & Y[8]) ^ S354;
    assign S356 = (X[4] & Y[7]) ^ S355;
    assign S357 = (X[5] & Y[6]) ^ S356;
    assign S358 = (X[6] & Y[5]) ^ S357;
    assign S359 = (X[7] & Y[4]) ^ S358;
    assign S360 = (X[8] & Y[3]) ^ S359;
    assign S361 = (X[9] & Y[2]) ^ S360;
    assign S362 = (X[10] & Y[1]) ^ S361;
    assign S363 = (X[11] & Y[0]) ^ S362;
    assign ClmulResult[11] = S363;
    assign S384 = X[0] & Y[12];
    assign S385 = (X[1] & Y[11]) ^ S384;
    assign S386 = (X[2] & Y[10]) ^ S385;
    assign S387 = (X[3] & Y[9]) ^ S386;
    assign S388 = (X[4] & Y[8]) ^ S387;
    assign S389 = (X[5] & Y[7]) ^ S388;
    assign S390 = (X[6] & Y[6]) ^ S389;
    assign S391 = (X[7] & Y[5]) ^ S390;
    assign S392 = (X[8] & Y[4]) ^ S391;
    assign S393 = (X[9] & Y[3]) ^ S392;
    assign S394 = (X[10] & Y[2]) ^ S393;
    assign S395 = (X[11] & Y[1]) ^ S394;
    assign S396 = (X[12] & Y[0]) ^ S395;
    assign ClmulResult[12] = S396;
    assign S416 = X[0] & Y[13];
    assign S417 = (X[1] & Y[12]) ^ S416;
    assign S418 = (X[2] & Y[11]) ^ S417;
    assign S419 = (X[3] & Y[10]) ^ S418;
    assign S420 = (X[4] & Y[9]) ^ S419;
    assign S421 = (X[5] & Y[8]) ^ S420;
    assign S422 = (X[6] & Y[7]) ^ S421;
    assign S423 = (X[7] & Y[6]) ^ S422;
    assign S424 = (X[8] & Y[5]) ^ S423;
    assign S425 = (X[9] & Y[4]) ^ S424;
    assign S426 = (X[10] & Y[3]) ^ S425;
    assign S427 = (X[11] & Y[2]) ^ S426;
    assign S428 = (X[12] & Y[1]) ^ S427;
    assign S429 = (X[13] & Y[0]) ^ S428;
    assign ClmulResult[13] = S429;
    assign S448 = X[0] & Y[14];
    assign S449 = (X[1] & Y[13]) ^ S448;
    assign S450 = (X[2] & Y[12]) ^ S449;
    assign S451 = (X[3] & Y[11]) ^ S450;
    assign S452 = (X[4] & Y[10]) ^ S451;
    assign S453 = (X[5] & Y[9]) ^ S452;
    assign S454 = (X[6] & Y[8]) ^ S453;
    assign S455 = (X[7] & Y[7]) ^ S454;
    assign S456 = (X[8] & Y[6]) ^ S455;
    assign S457 = (X[9] & Y[5]) ^ S456;
    assign S458 = (X[10] & Y[4]) ^ S457;
    assign S459 = (X[11] & Y[3]) ^ S458;
    assign S460 = (X[12] & Y[2]) ^ S459;
    assign S461 = (X[13] & Y[1]) ^ S460;
    assign S462 = (X[14] & Y[0]) ^ S461;
    assign ClmulResult[14] = S462;
    assign S480 = X[0] & Y[15];
    assign S481 = (X[1] & Y[14]) ^ S480;
    assign S482 = (X[2] & Y[13]) ^ S481;
    assign S483 = (X[3] & Y[12]) ^ S482;
    assign S484 = (X[4] & Y[11]) ^ S483;
    assign S485 = (X[5] & Y[10]) ^ S484;
    assign S486 = (X[6] & Y[9]) ^ S485;
    assign S487 = (X[7] & Y[8]) ^ S486;
    assign S488 = (X[8] & Y[7]) ^ S487;
    assign S489 = (X[9] & Y[6]) ^ S488;
    assign S490 = (X[10] & Y[5]) ^ S489;
    assign S491 = (X[11] & Y[4]) ^ S490;
    assign S492 = (X[12] & Y[3]) ^ S491;
    assign S493 = (X[13] & Y[2]) ^ S492;
    assign S494 = (X[14] & Y[1]) ^ S493;
    assign S495 = (X[15] & Y[0]) ^ S494;
    assign ClmulResult[15] = S495;
    assign S512 = X[0] & Y[16];
    assign S513 = (X[1] & Y[15]) ^ S512;
    assign S514 = (X[2] & Y[14]) ^ S513;
    assign S515 = (X[3] & Y[13]) ^ S514;
    assign S516 = (X[4] & Y[12]) ^ S515;
    assign S517 = (X[5] & Y[11]) ^ S516;
    assign S518 = (X[6] & Y[10]) ^ S517;
    assign S519 = (X[7] & Y[9]) ^ S518;
    assign S520 = (X[8] & Y[8]) ^ S519;
    assign S521 = (X[9] & Y[7]) ^ S520;
    assign S522 = (X[10] & Y[6]) ^ S521;
    assign S523 = (X[11] & Y[5]) ^ S522;
    assign S524 = (X[12] & Y[4]) ^ S523;
    assign S525 = (X[13] & Y[3]) ^ S524;
    assign S526 = (X[14] & Y[2]) ^ S525;
    assign S527 = (X[15] & Y[1]) ^ S526;
    assign S528 = (X[16] & Y[0]) ^ S527;
    assign ClmulResult[16] = S528;
    assign S544 = X[0] & Y[17];
    assign S545 = (X[1] & Y[16]) ^ S544;
    assign S546 = (X[2] & Y[15]) ^ S545;
    assign S547 = (X[3] & Y[14]) ^ S546;
    assign S548 = (X[4] & Y[13]) ^ S547;
    assign S549 = (X[5] & Y[12]) ^ S548;
    assign S550 = (X[6] & Y[11]) ^ S549;
    assign S551 = (X[7] & Y[10]) ^ S550;
    assign S552 = (X[8] & Y[9]) ^ S551;
    assign S553 = (X[9] & Y[8]) ^ S552;
    assign S554 = (X[10] & Y[7]) ^ S553;
    assign S555 = (X[11] & Y[6]) ^ S554;
    assign S556 = (X[12] & Y[5]) ^ S555;
    assign S557 = (X[13] & Y[4]) ^ S556;
    assign S558 = (X[14] & Y[3]) ^ S557;
    assign S559 = (X[15] & Y[2]) ^ S558;
    assign S560 = (X[16] & Y[1]) ^ S559;
    assign S561 = (X[17] & Y[0]) ^ S560;
    assign ClmulResult[17] = S561;
    assign S576 = X[0] & Y[18];
    assign S577 = (X[1] & Y[17]) ^ S576;
    assign S578 = (X[2] & Y[16]) ^ S577;
    assign S579 = (X[3] & Y[15]) ^ S578;
    assign S580 = (X[4] & Y[14]) ^ S579;
    assign S581 = (X[5] & Y[13]) ^ S580;
    assign S582 = (X[6] & Y[12]) ^ S581;
    assign S583 = (X[7] & Y[11]) ^ S582;
    assign S584 = (X[8] & Y[10]) ^ S583;
    assign S585 = (X[9] & Y[9]) ^ S584;
    assign S586 = (X[10] & Y[8]) ^ S585;
    assign S587 = (X[11] & Y[7]) ^ S586;
    assign S588 = (X[12] & Y[6]) ^ S587;
    assign S589 = (X[13] & Y[5]) ^ S588;
    assign S590 = (X[14] & Y[4]) ^ S589;
    assign S591 = (X[15] & Y[3]) ^ S590;
    assign S592 = (X[16] & Y[2]) ^ S591;
    assign S593 = (X[17] & Y[1]) ^ S592;
    assign S594 = (X[18] & Y[0]) ^ S593;
    assign ClmulResult[18] = S594;
    assign S608 = X[0] & Y[19];
    assign S609 = (X[1] & Y[18]) ^ S608;
    assign S610 = (X[2] & Y[17]) ^ S609;
    assign S611 = (X[3] & Y[16]) ^ S610;
    assign S612 = (X[4] & Y[15]) ^ S611;
    assign S613 = (X[5] & Y[14]) ^ S612;
    assign S614 = (X[6] & Y[13]) ^ S613;
    assign S615 = (X[7] & Y[12]) ^ S614;
    assign S616 = (X[8] & Y[11]) ^ S615;
    assign S617 = (X[9] & Y[10]) ^ S616;
    assign S618 = (X[10] & Y[9]) ^ S617;
    assign S619 = (X[11] & Y[8]) ^ S618;
    assign S620 = (X[12] & Y[7]) ^ S619;
    assign S621 = (X[13] & Y[6]) ^ S620;
    assign S622 = (X[14] & Y[5]) ^ S621;
    assign S623 = (X[15] & Y[4]) ^ S622;
    assign S624 = (X[16] & Y[3]) ^ S623;
    assign S625 = (X[17] & Y[2]) ^ S624;
    assign S626 = (X[18] & Y[1]) ^ S625;
    assign S627 = (X[19] & Y[0]) ^ S626;
    assign ClmulResult[19] = S627;
    assign S640 = X[0] & Y[20];
    assign S641 = (X[1] & Y[19]) ^ S640;
    assign S642 = (X[2] & Y[18]) ^ S641;
    assign S643 = (X[3] & Y[17]) ^ S642;
    assign S644 = (X[4] & Y[16]) ^ S643;
    assign S645 = (X[5] & Y[15]) ^ S644;
    assign S646 = (X[6] & Y[14]) ^ S645;
    assign S647 = (X[7] & Y[13]) ^ S646;
    assign S648 = (X[8] & Y[12]) ^ S647;
    assign S649 = (X[9] & Y[11]) ^ S648;
    assign S650 = (X[10] & Y[10]) ^ S649;
    assign S651 = (X[11] & Y[9]) ^ S650;
    assign S652 = (X[12] & Y[8]) ^ S651;
    assign S653 = (X[13] & Y[7]) ^ S652;
    assign S654 = (X[14] & Y[6]) ^ S653;
    assign S655 = (X[15] & Y[5]) ^ S654;
    assign S656 = (X[16] & Y[4]) ^ S655;
    assign S657 = (X[17] & Y[3]) ^ S656;
    assign S658 = (X[18] & Y[2]) ^ S657;
    assign S659 = (X[19] & Y[1]) ^ S658;
    assign S660 = (X[20] & Y[0]) ^ S659;
    assign ClmulResult[20] = S660;
    assign S672 = X[0] & Y[21];
    assign S673 = (X[1] & Y[20]) ^ S672;
    assign S674 = (X[2] & Y[19]) ^ S673;
    assign S675 = (X[3] & Y[18]) ^ S674;
    assign S676 = (X[4] & Y[17]) ^ S675;
    assign S677 = (X[5] & Y[16]) ^ S676;
    assign S678 = (X[6] & Y[15]) ^ S677;
    assign S679 = (X[7] & Y[14]) ^ S678;
    assign S680 = (X[8] & Y[13]) ^ S679;
    assign S681 = (X[9] & Y[12]) ^ S680;
    assign S682 = (X[10] & Y[11]) ^ S681;
    assign S683 = (X[11] & Y[10]) ^ S682;
    assign S684 = (X[12] & Y[9]) ^ S683;
    assign S685 = (X[13] & Y[8]) ^ S684;
    assign S686 = (X[14] & Y[7]) ^ S685;
    assign S687 = (X[15] & Y[6]) ^ S686;
    assign S688 = (X[16] & Y[5]) ^ S687;
    assign S689 = (X[17] & Y[4]) ^ S688;
    assign S690 = (X[18] & Y[3]) ^ S689;
    assign S691 = (X[19] & Y[2]) ^ S690;
    assign S692 = (X[20] & Y[1]) ^ S691;
    assign S693 = (X[21] & Y[0]) ^ S692;
    assign ClmulResult[21] = S693;
    assign S704 = X[0] & Y[22];
    assign S705 = (X[1] & Y[21]) ^ S704;
    assign S706 = (X[2] & Y[20]) ^ S705;
    assign S707 = (X[3] & Y[19]) ^ S706;
    assign S708 = (X[4] & Y[18]) ^ S707;
    assign S709 = (X[5] & Y[17]) ^ S708;
    assign S710 = (X[6] & Y[16]) ^ S709;
    assign S711 = (X[7] & Y[15]) ^ S710;
    assign S712 = (X[8] & Y[14]) ^ S711;
    assign S713 = (X[9] & Y[13]) ^ S712;
    assign S714 = (X[10] & Y[12]) ^ S713;
    assign S715 = (X[11] & Y[11]) ^ S714;
    assign S716 = (X[12] & Y[10]) ^ S715;
    assign S717 = (X[13] & Y[9]) ^ S716;
    assign S718 = (X[14] & Y[8]) ^ S717;
    assign S719 = (X[15] & Y[7]) ^ S718;
    assign S720 = (X[16] & Y[6]) ^ S719;
    assign S721 = (X[17] & Y[5]) ^ S720;
    assign S722 = (X[18] & Y[4]) ^ S721;
    assign S723 = (X[19] & Y[3]) ^ S722;
    assign S724 = (X[20] & Y[2]) ^ S723;
    assign S725 = (X[21] & Y[1]) ^ S724;
    assign S726 = (X[22] & Y[0]) ^ S725;
    assign ClmulResult[22] = S726;
    assign S736 = X[0] & Y[23];
    assign S737 = (X[1] & Y[22]) ^ S736;
    assign S738 = (X[2] & Y[21]) ^ S737;
    assign S739 = (X[3] & Y[20]) ^ S738;
    assign S740 = (X[4] & Y[19]) ^ S739;
    assign S741 = (X[5] & Y[18]) ^ S740;
    assign S742 = (X[6] & Y[17]) ^ S741;
    assign S743 = (X[7] & Y[16]) ^ S742;
    assign S744 = (X[8] & Y[15]) ^ S743;
    assign S745 = (X[9] & Y[14]) ^ S744;
    assign S746 = (X[10] & Y[13]) ^ S745;
    assign S747 = (X[11] & Y[12]) ^ S746;
    assign S748 = (X[12] & Y[11]) ^ S747;
    assign S749 = (X[13] & Y[10]) ^ S748;
    assign S750 = (X[14] & Y[9]) ^ S749;
    assign S751 = (X[15] & Y[8]) ^ S750;
    assign S752 = (X[16] & Y[7]) ^ S751;
    assign S753 = (X[17] & Y[6]) ^ S752;
    assign S754 = (X[18] & Y[5]) ^ S753;
    assign S755 = (X[19] & Y[4]) ^ S754;
    assign S756 = (X[20] & Y[3]) ^ S755;
    assign S757 = (X[21] & Y[2]) ^ S756;
    assign S758 = (X[22] & Y[1]) ^ S757;
    assign S759 = (X[23] & Y[0]) ^ S758;
    assign ClmulResult[23] = S759;
    assign S768 = X[0] & Y[24];
    assign S769 = (X[1] & Y[23]) ^ S768;
    assign S770 = (X[2] & Y[22]) ^ S769;
    assign S771 = (X[3] & Y[21]) ^ S770;
    assign S772 = (X[4] & Y[20]) ^ S771;
    assign S773 = (X[5] & Y[19]) ^ S772;
    assign S774 = (X[6] & Y[18]) ^ S773;
    assign S775 = (X[7] & Y[17]) ^ S774;
    assign S776 = (X[8] & Y[16]) ^ S775;
    assign S777 = (X[9] & Y[15]) ^ S776;
    assign S778 = (X[10] & Y[14]) ^ S777;
    assign S779 = (X[11] & Y[13]) ^ S778;
    assign S780 = (X[12] & Y[12]) ^ S779;
    assign S781 = (X[13] & Y[11]) ^ S780;
    assign S782 = (X[14] & Y[10]) ^ S781;
    assign S783 = (X[15] & Y[9]) ^ S782;
    assign S784 = (X[16] & Y[8]) ^ S783;
    assign S785 = (X[17] & Y[7]) ^ S784;
    assign S786 = (X[18] & Y[6]) ^ S785;
    assign S787 = (X[19] & Y[5]) ^ S786;
    assign S788 = (X[20] & Y[4]) ^ S787;
    assign S789 = (X[21] & Y[3]) ^ S788;
    assign S790 = (X[22] & Y[2]) ^ S789;
    assign S791 = (X[23] & Y[1]) ^ S790;
    assign S792 = (X[24] & Y[0]) ^ S791;
    assign ClmulResult[24] = S792;
    assign S800 = X[0] & Y[25];
    assign S801 = (X[1] & Y[24]) ^ S800;
    assign S802 = (X[2] & Y[23]) ^ S801;
    assign S803 = (X[3] & Y[22]) ^ S802;
    assign S804 = (X[4] & Y[21]) ^ S803;
    assign S805 = (X[5] & Y[20]) ^ S804;
    assign S806 = (X[6] & Y[19]) ^ S805;
    assign S807 = (X[7] & Y[18]) ^ S806;
    assign S808 = (X[8] & Y[17]) ^ S807;
    assign S809 = (X[9] & Y[16]) ^ S808;
    assign S810 = (X[10] & Y[15]) ^ S809;
    assign S811 = (X[11] & Y[14]) ^ S810;
    assign S812 = (X[12] & Y[13]) ^ S811;
    assign S813 = (X[13] & Y[12]) ^ S812;
    assign S814 = (X[14] & Y[11]) ^ S813;
    assign S815 = (X[15] & Y[10]) ^ S814;
    assign S816 = (X[16] & Y[9]) ^ S815;
    assign S817 = (X[17] & Y[8]) ^ S816;
    assign S818 = (X[18] & Y[7]) ^ S817;
    assign S819 = (X[19] & Y[6]) ^ S818;
    assign S820 = (X[20] & Y[5]) ^ S819;
    assign S821 = (X[21] & Y[4]) ^ S820;
    assign S822 = (X[22] & Y[3]) ^ S821;
    assign S823 = (X[23] & Y[2]) ^ S822;
    assign S824 = (X[24] & Y[1]) ^ S823;
    assign S825 = (X[25] & Y[0]) ^ S824;
    assign ClmulResult[25] = S825;
    assign S832 = X[0] & Y[26];
    assign S833 = (X[1] & Y[25]) ^ S832;
    assign S834 = (X[2] & Y[24]) ^ S833;
    assign S835 = (X[3] & Y[23]) ^ S834;
    assign S836 = (X[4] & Y[22]) ^ S835;
    assign S837 = (X[5] & Y[21]) ^ S836;
    assign S838 = (X[6] & Y[20]) ^ S837;
    assign S839 = (X[7] & Y[19]) ^ S838;
    assign S840 = (X[8] & Y[18]) ^ S839;
    assign S841 = (X[9] & Y[17]) ^ S840;
    assign S842 = (X[10] & Y[16]) ^ S841;
    assign S843 = (X[11] & Y[15]) ^ S842;
    assign S844 = (X[12] & Y[14]) ^ S843;
    assign S845 = (X[13] & Y[13]) ^ S844;
    assign S846 = (X[14] & Y[12]) ^ S845;
    assign S847 = (X[15] & Y[11]) ^ S846;
    assign S848 = (X[16] & Y[10]) ^ S847;
    assign S849 = (X[17] & Y[9]) ^ S848;
    assign S850 = (X[18] & Y[8]) ^ S849;
    assign S851 = (X[19] & Y[7]) ^ S850;
    assign S852 = (X[20] & Y[6]) ^ S851;
    assign S853 = (X[21] & Y[5]) ^ S852;
    assign S854 = (X[22] & Y[4]) ^ S853;
    assign S855 = (X[23] & Y[3]) ^ S854;
    assign S856 = (X[24] & Y[2]) ^ S855;
    assign S857 = (X[25] & Y[1]) ^ S856;
    assign S858 = (X[26] & Y[0]) ^ S857;
    assign ClmulResult[26] = S858;
    assign S864 = X[0] & Y[27];
    assign S865 = (X[1] & Y[26]) ^ S864;
    assign S866 = (X[2] & Y[25]) ^ S865;
    assign S867 = (X[3] & Y[24]) ^ S866;
    assign S868 = (X[4] & Y[23]) ^ S867;
    assign S869 = (X[5] & Y[22]) ^ S868;
    assign S870 = (X[6] & Y[21]) ^ S869;
    assign S871 = (X[7] & Y[20]) ^ S870;
    assign S872 = (X[8] & Y[19]) ^ S871;
    assign S873 = (X[9] & Y[18]) ^ S872;
    assign S874 = (X[10] & Y[17]) ^ S873;
    assign S875 = (X[11] & Y[16]) ^ S874;
    assign S876 = (X[12] & Y[15]) ^ S875;
    assign S877 = (X[13] & Y[14]) ^ S876;
    assign S878 = (X[14] & Y[13]) ^ S877;
    assign S879 = (X[15] & Y[12]) ^ S878;
    assign S880 = (X[16] & Y[11]) ^ S879;
    assign S881 = (X[17] & Y[10]) ^ S880;
    assign S882 = (X[18] & Y[9]) ^ S881;
    assign S883 = (X[19] & Y[8]) ^ S882;
    assign S884 = (X[20] & Y[7]) ^ S883;
    assign S885 = (X[21] & Y[6]) ^ S884;
    assign S886 = (X[22] & Y[5]) ^ S885;
    assign S887 = (X[23] & Y[4]) ^ S886;
    assign S888 = (X[24] & Y[3]) ^ S887;
    assign S889 = (X[25] & Y[2]) ^ S888;
    assign S890 = (X[26] & Y[1]) ^ S889;
    assign S891 = (X[27] & Y[0]) ^ S890;
    assign ClmulResult[27] = S891;
    assign S896 = X[0] & Y[28];
    assign S897 = (X[1] & Y[27]) ^ S896;
    assign S898 = (X[2] & Y[26]) ^ S897;
    assign S899 = (X[3] & Y[25]) ^ S898;
    assign S900 = (X[4] & Y[24]) ^ S899;
    assign S901 = (X[5] & Y[23]) ^ S900;
    assign S902 = (X[6] & Y[22]) ^ S901;
    assign S903 = (X[7] & Y[21]) ^ S902;
    assign S904 = (X[8] & Y[20]) ^ S903;
    assign S905 = (X[9] & Y[19]) ^ S904;
    assign S906 = (X[10] & Y[18]) ^ S905;
    assign S907 = (X[11] & Y[17]) ^ S906;
    assign S908 = (X[12] & Y[16]) ^ S907;
    assign S909 = (X[13] & Y[15]) ^ S908;
    assign S910 = (X[14] & Y[14]) ^ S909;
    assign S911 = (X[15] & Y[13]) ^ S910;
    assign S912 = (X[16] & Y[12]) ^ S911;
    assign S913 = (X[17] & Y[11]) ^ S912;
    assign S914 = (X[18] & Y[10]) ^ S913;
    assign S915 = (X[19] & Y[9]) ^ S914;
    assign S916 = (X[20] & Y[8]) ^ S915;
    assign S917 = (X[21] & Y[7]) ^ S916;
    assign S918 = (X[22] & Y[6]) ^ S917;
    assign S919 = (X[23] & Y[5]) ^ S918;
    assign S920 = (X[24] & Y[4]) ^ S919;
    assign S921 = (X[25] & Y[3]) ^ S920;
    assign S922 = (X[26] & Y[2]) ^ S921;
    assign S923 = (X[27] & Y[1]) ^ S922;
    assign S924 = (X[28] & Y[0]) ^ S923;
    assign ClmulResult[28] = S924;
    assign S928 = X[0] & Y[29];
    assign S929 = (X[1] & Y[28]) ^ S928;
    assign S930 = (X[2] & Y[27]) ^ S929;
    assign S931 = (X[3] & Y[26]) ^ S930;
    assign S932 = (X[4] & Y[25]) ^ S931;
    assign S933 = (X[5] & Y[24]) ^ S932;
    assign S934 = (X[6] & Y[23]) ^ S933;
    assign S935 = (X[7] & Y[22]) ^ S934;
    assign S936 = (X[8] & Y[21]) ^ S935;
    assign S937 = (X[9] & Y[20]) ^ S936;
    assign S938 = (X[10] & Y[19]) ^ S937;
    assign S939 = (X[11] & Y[18]) ^ S938;
    assign S940 = (X[12] & Y[17]) ^ S939;
    assign S941 = (X[13] & Y[16]) ^ S940;
    assign S942 = (X[14] & Y[15]) ^ S941;
    assign S943 = (X[15] & Y[14]) ^ S942;
    assign S944 = (X[16] & Y[13]) ^ S943;
    assign S945 = (X[17] & Y[12]) ^ S944;
    assign S946 = (X[18] & Y[11]) ^ S945;
    assign S947 = (X[19] & Y[10]) ^ S946;
    assign S948 = (X[20] & Y[9]) ^ S947;
    assign S949 = (X[21] & Y[8]) ^ S948;
    assign S950 = (X[22] & Y[7]) ^ S949;
    assign S951 = (X[23] & Y[6]) ^ S950;
    assign S952 = (X[24] & Y[5]) ^ S951;
    assign S953 = (X[25] & Y[4]) ^ S952;
    assign S954 = (X[26] & Y[3]) ^ S953;
    assign S955 = (X[27] & Y[2]) ^ S954;
    assign S956 = (X[28] & Y[1]) ^ S955;
    assign S957 = (X[29] & Y[0]) ^ S956;
    assign ClmulResult[29] = S957;
    assign S960 = X[0] & Y[30];
    assign S961 = (X[1] & Y[29]) ^ S960;
    assign S962 = (X[2] & Y[28]) ^ S961;
    assign S963 = (X[3] & Y[27]) ^ S962;
    assign S964 = (X[4] & Y[26]) ^ S963;
    assign S965 = (X[5] & Y[25]) ^ S964;
    assign S966 = (X[6] & Y[24]) ^ S965;
    assign S967 = (X[7] & Y[23]) ^ S966;
    assign S968 = (X[8] & Y[22]) ^ S967;
    assign S969 = (X[9] & Y[21]) ^ S968;
    assign S970 = (X[10] & Y[20]) ^ S969;
    assign S971 = (X[11] & Y[19]) ^ S970;
    assign S972 = (X[12] & Y[18]) ^ S971;
    assign S973 = (X[13] & Y[17]) ^ S972;
    assign S974 = (X[14] & Y[16]) ^ S973;
    assign S975 = (X[15] & Y[15]) ^ S974;
    assign S976 = (X[16] & Y[14]) ^ S975;
    assign S977 = (X[17] & Y[13]) ^ S976;
    assign S978 = (X[18] & Y[12]) ^ S977;
    assign S979 = (X[19] & Y[11]) ^ S978;
    assign S980 = (X[20] & Y[10]) ^ S979;
    assign S981 = (X[21] & Y[9]) ^ S980;
    assign S982 = (X[22] & Y[8]) ^ S981;
    assign S983 = (X[23] & Y[7]) ^ S982;
    assign S984 = (X[24] & Y[6]) ^ S983;
    assign S985 = (X[25] & Y[5]) ^ S984;
    assign S986 = (X[26] & Y[4]) ^ S985;
    assign S987 = (X[27] & Y[3]) ^ S986;
    assign S988 = (X[28] & Y[2]) ^ S987;
    assign S989 = (X[29] & Y[1]) ^ S988;
    assign S990 = (X[30] & Y[0]) ^ S989;
    assign ClmulResult[30] = S990;
    assign S992 = X[0] & Y[31];
    assign S993 = (X[1] & Y[30]) ^ S992;
    assign S994 = (X[2] & Y[29]) ^ S993;
    assign S995 = (X[3] & Y[28]) ^ S994;
    assign S996 = (X[4] & Y[27]) ^ S995;
    assign S997 = (X[5] & Y[26]) ^ S996;
    assign S998 = (X[6] & Y[25]) ^ S997;
    assign S999 = (X[7] & Y[24]) ^ S998;
    assign S1000 = (X[8] & Y[23]) ^ S999;
    assign S1001 = (X[9] & Y[22]) ^ S1000;
    assign S1002 = (X[10] & Y[21]) ^ S1001;
    assign S1003 = (X[11] & Y[20]) ^ S1002;
    assign S1004 = (X[12] & Y[19]) ^ S1003;
    assign S1005 = (X[13] & Y[18]) ^ S1004;
    assign S1006 = (X[14] & Y[17]) ^ S1005;
    assign S1007 = (X[15] & Y[16]) ^ S1006;
    assign S1008 = (X[16] & Y[15]) ^ S1007;
    assign S1009 = (X[17] & Y[14]) ^ S1008;
    assign S1010 = (X[18] & Y[13]) ^ S1009;
    assign S1011 = (X[19] & Y[12]) ^ S1010;
    assign S1012 = (X[20] & Y[11]) ^ S1011;
    assign S1013 = (X[21] & Y[10]) ^ S1012;
    assign S1014 = (X[22] & Y[9]) ^ S1013;
    assign S1015 = (X[23] & Y[8]) ^ S1014;
    assign S1016 = (X[24] & Y[7]) ^ S1015;
    assign S1017 = (X[25] & Y[6]) ^ S1016;
    assign S1018 = (X[26] & Y[5]) ^ S1017;
    assign S1019 = (X[27] & Y[4]) ^ S1018;
    assign S1020 = (X[28] & Y[3]) ^ S1019;
    assign S1021 = (X[29] & Y[2]) ^ S1020;
    assign S1022 = (X[30] & Y[1]) ^ S1021;
    assign S1023 = (X[31] & Y[0]) ^ S1022;
    assign ClmulResult[31] = S1023;

  end
endmodule


