
///////////////////////////////////////////
// popccnt.sv
// Written: Kevin Kim <kekim@hmc.edu>
// Modified: 2/4/2023
//
// Purpose: Population Count
// 
// A component of the CORE-V-WALLY configurable RISC-V project.
// 
// Copyright (C) 2021-23 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

module popcntcsa2 #(parameter WIDTH = 16) (
  input logic  [WIDTH-1:0]            a,    // number to count total ones
  output logic [$clog2(WIDTH):0]  s  // the total number of ones
);
if (WIDTH == 8)begin

  assign {w0_0_7, w0_0_6, w0_0_5, w0_0_4, w0_0_3, w0_0_2, w0_0_1, w0_0_0} = a;
logic w1_0_0;
logic w0_1_15;
csan2 csan0_0_7_0_0_6_X_X_X(w0_0_7, w0_0_6, w1_0_0, w0_1_15);
logic w1_0_1;
logic w0_1_13;
csan2 csan0_0_5_0_0_4_X_X_X(w0_0_5, w0_0_4, w1_0_1, w0_1_13);
logic w1_0_2;
logic w0_1_11;
csan2 csan0_0_3_0_0_2_X_X_X(w0_0_3, w0_0_2, w1_0_2, w0_1_11);
logic w1_0_3;
logic w0_1_9;
csan2 csan0_0_1_0_0_0_X_X_X(w0_0_1, w0_0_0, w1_0_3, w0_1_9);
logic w1_0_4;
logic w0_2_23;
csan2 csan0_1_15_0_1_13_X_X_X(w0_1_15, w0_1_13, w1_0_4, w0_2_23);
logic w1_0_5;
logic w0_2_19;
csan2 csan0_1_11_0_1_9_X_X_X(w0_1_11, w0_1_9, w1_0_5, w0_2_19);
logic w1_0_6;
logic w0_3_31;
csan2 csan0_2_23_0_2_19_X_X_X(w0_2_23, w0_2_19, w1_0_6, w0_3_31);
assign s0 = w0_3_31;
logic w2_0_0;
logic w1_1_8;
csan2 csan1_0_0_1_0_1_X_X_X(w1_0_0, w1_0_1, w2_0_0, w1_1_8);
logic w2_0_1;
logic w1_1_10;
csan2 csan1_0_2_1_0_3_X_X_X(w1_0_2, w1_0_3, w2_0_1, w1_1_10);
logic w2_0_2;
logic w1_1_12;
csan2 csan1_0_4_1_0_5_X_X_X(w1_0_4, w1_0_5, w2_0_2, w1_1_12);
logic w2_0_3;
logic w1_2_14;
csan2 csan1_0_6_1_1_8_X_X_X(w1_0_6, w1_1_8, w2_0_3, w1_2_14);
logic w2_0_4;
logic w1_2_18;
csan2 csan1_1_10_1_1_12_X_X_X(w1_1_10, w1_1_12, w2_0_4, w1_2_18);
logic w2_0_5;
logic w1_3_22;
csan2 csan1_2_14_1_2_18_X_X_X(w1_2_14, w1_2_18, w2_0_5, w1_3_22);
assign s1 = w1_3_22;
logic w3_0_0;
logic w2_1_8;
csan2 csan2_0_0_2_0_1_X_X_X(w2_0_0, w2_0_1, w3_0_0, w2_1_8);
logic w3_0_1;
logic w2_1_10;
csan2 csan2_0_2_2_0_3_X_X_X(w2_0_2, w2_0_3, w3_0_1, w2_1_10);
logic w3_0_2;
logic w2_1_12;
csan2 csan2_0_4_2_0_5_X_X_X(w2_0_4, w2_0_5, w3_0_2, w2_1_12);
logic w3_0_3;
logic w2_2_16;
csan2 csan2_1_8_2_1_10_X_X_X(w2_1_8, w2_1_10, w3_0_3, w2_2_16);
logic w3_0_4;
logic w2_3_20;
csan2 csan2_1_12_2_2_16_X_X_X(w2_1_12, w2_2_16, w3_0_4, w2_3_20);
assign s2 = w2_3_20;
logic w4_0_0;
logic w3_1_8;
csan2 csan3_0_0_3_0_1_X_X_X(w3_0_0, w3_0_1, w4_0_0, w3_1_8);
logic w4_0_1;
logic w3_1_10;
csan2 csan3_0_2_3_0_3_X_X_X(w3_0_2, w3_0_3, w4_0_1, w3_1_10);
logic w4_0_2;
logic w3_2_12;
csan2 csan3_0_4_3_1_8_X_X_X(w3_0_4, w3_1_8, w4_0_2, w3_2_12);
logic w4_0_3;
logic w3_3_18;
csan2 csan3_1_10_3_2_12_X_X_X(w3_1_10, w3_2_12, w4_0_3, w3_3_18);
assign s3 = w3_3_18;
  assign s = {s3,s2,s1,s0};
end
else if (WIDTH == 16) begin
  assign {w0_0_15, w0_0_14, w0_0_13, w0_0_12, w0_0_11, w0_0_10, w0_0_9, w0_0_8, w0_0_7, w0_0_6, w0_0_5, w0_0_4, w0_0_3, w0_0_2, w0_0_1, w0_0_0} = a;
  logic w1_0_0;
  logic w0_1_31;
  csan2 csan0_0_15_0_0_14_X_X_X(w0_0_15, w0_0_14, w1_0_0, w0_1_31);
  logic w1_0_1;
  logic w0_1_29;
  csan2 csan0_0_13_0_0_12_X_X_X(w0_0_13, w0_0_12, w1_0_1, w0_1_29);
  logic w1_0_2;
  logic w0_1_27;
  csan2 csan0_0_11_0_0_10_X_X_X(w0_0_11, w0_0_10, w1_0_2, w0_1_27);
  logic w1_0_3;
  logic w0_1_25;
  csan2 csan0_0_9_0_0_8_X_X_X(w0_0_9, w0_0_8, w1_0_3, w0_1_25);
  logic w1_0_4;
  logic w0_1_23;
  csan2 csan0_0_7_0_0_6_X_X_X(w0_0_7, w0_0_6, w1_0_4, w0_1_23);
  logic w1_0_5;
  logic w0_1_21;
  csan2 csan0_0_5_0_0_4_X_X_X(w0_0_5, w0_0_4, w1_0_5, w0_1_21);
  logic w1_0_6;
  logic w0_1_19;
  csan2 csan0_0_3_0_0_2_X_X_X(w0_0_3, w0_0_2, w1_0_6, w0_1_19);
  logic w1_0_7;
  logic w0_1_17;
  csan2 csan0_0_1_0_0_0_X_X_X(w0_0_1, w0_0_0, w1_0_7, w0_1_17);
  logic w1_0_8;
  logic w0_2_47;
  csan2 csan0_1_31_0_1_29_X_X_X(w0_1_31, w0_1_29, w1_0_8, w0_2_47);
  logic w1_0_9;
  logic w0_2_43;
  csan2 csan0_1_27_0_1_25_X_X_X(w0_1_27, w0_1_25, w1_0_9, w0_2_43);
  logic w1_0_10;
  logic w0_2_39;
  csan2 csan0_1_23_0_1_21_X_X_X(w0_1_23, w0_1_21, w1_0_10, w0_2_39);
  logic w1_0_11;
  logic w0_2_35;
  csan2 csan0_1_19_0_1_17_X_X_X(w0_1_19, w0_1_17, w1_0_11, w0_2_35);
  logic w1_0_12;
  logic w0_3_63;
  csan2 csan0_2_47_0_2_43_X_X_X(w0_2_47, w0_2_43, w1_0_12, w0_3_63);
  logic w1_0_13;
  logic w0_3_55;
  csan2 csan0_2_39_0_2_35_X_X_X(w0_2_39, w0_2_35, w1_0_13, w0_3_55);
  logic w1_0_14;
  logic w0_4_79;
  csan2 csan0_3_63_0_3_55_X_X_X(w0_3_63, w0_3_55, w1_0_14, w0_4_79);
  assign s0 = w0_4_79;
  logic w2_0_0;
  logic w1_1_16;
  csan2 csan1_0_0_1_0_1_X_X_X(w1_0_0, w1_0_1, w2_0_0, w1_1_16);
  logic w2_0_1;
  logic w1_1_18;
  csan2 csan1_0_2_1_0_3_X_X_X(w1_0_2, w1_0_3, w2_0_1, w1_1_18);
  logic w2_0_2;
  logic w1_1_20;
  csan2 csan1_0_4_1_0_5_X_X_X(w1_0_4, w1_0_5, w2_0_2, w1_1_20);
  logic w2_0_3;
  logic w1_1_22;
  csan2 csan1_0_6_1_0_7_X_X_X(w1_0_6, w1_0_7, w2_0_3, w1_1_22);
  logic w2_0_4;
  logic w1_1_24;
  csan2 csan1_0_8_1_0_9_X_X_X(w1_0_8, w1_0_9, w2_0_4, w1_1_24);
  logic w2_0_5;
  logic w1_1_26;
  csan2 csan1_0_10_1_0_11_X_X_X(w1_0_10, w1_0_11, w2_0_5, w1_1_26);
  logic w2_0_6;
  logic w1_1_28;
  csan2 csan1_0_12_1_0_13_X_X_X(w1_0_12, w1_0_13, w2_0_6, w1_1_28);
  logic w2_0_7;
  logic w1_2_30;
  csan2 csan1_0_14_1_1_16_X_X_X(w1_0_14, w1_1_16, w2_0_7, w1_2_30);
  logic w2_0_8;
  logic w1_2_34;
  csan2 csan1_1_18_1_1_20_X_X_X(w1_1_18, w1_1_20, w2_0_8, w1_2_34);
  logic w2_0_9;
  logic w1_2_38;
  csan2 csan1_1_22_1_1_24_X_X_X(w1_1_22, w1_1_24, w2_0_9, w1_2_38);
  logic w2_0_10;
  logic w1_2_42;
  csan2 csan1_1_26_1_1_28_X_X_X(w1_1_26, w1_1_28, w2_0_10, w1_2_42);
  logic w2_0_11;
  logic w1_3_46;
  csan2 csan1_2_30_1_2_34_X_X_X(w1_2_30, w1_2_34, w2_0_11, w1_3_46);
  logic w2_0_12;
  logic w1_3_54;
  csan2 csan1_2_38_1_2_42_X_X_X(w1_2_38, w1_2_42, w2_0_12, w1_3_54);
  logic w2_0_13;
  logic w1_4_62;
  csan2 csan1_3_46_1_3_54_X_X_X(w1_3_46, w1_3_54, w2_0_13, w1_4_62);
  assign s1 = w1_4_62;
  logic w3_0_0;
  logic w2_1_16;
  csan2 csan2_0_0_2_0_1_X_X_X(w2_0_0, w2_0_1, w3_0_0, w2_1_16);
  logic w3_0_1;
  logic w2_1_18;
  csan2 csan2_0_2_2_0_3_X_X_X(w2_0_2, w2_0_3, w3_0_1, w2_1_18);
  logic w3_0_2;
  logic w2_1_20;
  csan2 csan2_0_4_2_0_5_X_X_X(w2_0_4, w2_0_5, w3_0_2, w2_1_20);
  logic w3_0_3;
  logic w2_1_22;
  csan2 csan2_0_6_2_0_7_X_X_X(w2_0_6, w2_0_7, w3_0_3, w2_1_22);
  logic w3_0_4;
  logic w2_1_24;
  csan2 csan2_0_8_2_0_9_X_X_X(w2_0_8, w2_0_9, w3_0_4, w2_1_24);
  logic w3_0_5;
  logic w2_1_26;
  csan2 csan2_0_10_2_0_11_X_X_X(w2_0_10, w2_0_11, w3_0_5, w2_1_26);
  logic w3_0_6;
  logic w2_1_28;
  csan2 csan2_0_12_2_0_13_X_X_X(w2_0_12, w2_0_13, w3_0_6, w2_1_28);
  logic w3_0_7;
  logic w2_2_32;
  csan2 csan2_1_16_2_1_18_X_X_X(w2_1_16, w2_1_18, w3_0_7, w2_2_32);
  logic w3_0_8;
  logic w2_2_36;
  csan2 csan2_1_20_2_1_22_X_X_X(w2_1_20, w2_1_22, w3_0_8, w2_2_36);
  logic w3_0_9;
  logic w2_2_40;
  csan2 csan2_1_24_2_1_26_X_X_X(w2_1_24, w2_1_26, w3_0_9, w2_2_40);
  logic w3_0_10;
  logic w2_3_44;
  csan2 csan2_1_28_2_2_32_X_X_X(w2_1_28, w2_2_32, w3_0_10, w2_3_44);
  logic w3_0_11;
  logic w2_3_52;
  csan2 csan2_2_36_2_2_40_X_X_X(w2_2_36, w2_2_40, w3_0_11, w2_3_52);
  logic w3_0_12;
  logic w2_4_60;
  csan2 csan2_3_44_2_3_52_X_X_X(w2_3_44, w2_3_52, w3_0_12, w2_4_60);
  assign s2 = w2_4_60;
  logic w4_0_0;
  logic w3_1_16;
  csan2 csan3_0_0_3_0_1_X_X_X(w3_0_0, w3_0_1, w4_0_0, w3_1_16);
  logic w4_0_1;
  logic w3_1_18;
  csan2 csan3_0_2_3_0_3_X_X_X(w3_0_2, w3_0_3, w4_0_1, w3_1_18);
  logic w4_0_2;
  logic w3_1_20;
  csan2 csan3_0_4_3_0_5_X_X_X(w3_0_4, w3_0_5, w4_0_2, w3_1_20);
  logic w4_0_3;
  logic w3_1_22;
  csan2 csan3_0_6_3_0_7_X_X_X(w3_0_6, w3_0_7, w4_0_3, w3_1_22);
  logic w4_0_4;
  logic w3_1_24;
  csan2 csan3_0_8_3_0_9_X_X_X(w3_0_8, w3_0_9, w4_0_4, w3_1_24);
  logic w4_0_5;
  logic w3_1_26;
  csan2 csan3_0_10_3_0_11_X_X_X(w3_0_10, w3_0_11, w4_0_5, w3_1_26);
  logic w4_0_6;
  logic w3_2_28;
  csan2 csan3_0_12_3_1_16_X_X_X(w3_0_12, w3_1_16, w4_0_6, w3_2_28);
  logic w4_0_7;
  logic w3_2_34;
  csan2 csan3_1_18_3_1_20_X_X_X(w3_1_18, w3_1_20, w4_0_7, w3_2_34);
  logic w4_0_8;
  logic w3_2_38;
  csan2 csan3_1_22_3_1_24_X_X_X(w3_1_22, w3_1_24, w4_0_8, w3_2_38);
  logic w4_0_9;
  logic w3_3_42;
  csan2 csan3_1_26_3_2_28_X_X_X(w3_1_26, w3_2_28, w4_0_9, w3_3_42);
  logic w4_0_10;
  logic w3_3_50;
  csan2 csan3_2_34_3_2_38_X_X_X(w3_2_34, w3_2_38, w4_0_10, w3_3_50);
  logic w4_0_11;
  logic w3_4_58;
  csan2 csan3_3_42_3_3_50_X_X_X(w3_3_42, w3_3_50, w4_0_11, w3_4_58);
  assign s3 = w3_4_58;
  logic w5_0_0;
  logic w4_1_16;
  csan1 csan4_0_0_4_0_1_X_X_X(w4_0_0, w4_0_1, w4_1_16);
  logic w5_0_1;
  logic w4_1_18;
  csan1 csan4_0_2_4_0_3_X_X_X(w4_0_2, w4_0_3, w4_1_18);
  logic w5_0_2;
  logic w4_1_20;
  csan1 csan4_0_4_4_0_5_X_X_X(w4_0_4, w4_0_5, w4_1_20);
  logic w5_0_3;
  logic w4_1_22;
  csan1 csan4_0_6_4_0_7_X_X_X(w4_0_6, w4_0_7, w4_1_22);
  logic w5_0_4;
  logic w4_1_24;
  csan1 csan4_0_8_4_0_9_X_X_X(w4_0_8, w4_0_9, w4_1_24);
  logic w5_0_5;
  logic w4_1_26;
  csan1 csan4_0_10_4_0_11_X_X_X(w4_0_10, w4_0_11, w4_1_26);
  logic w5_0_6;
  logic w4_2_32;
  csan1 csan4_1_16_4_1_18_X_X_X(w4_1_16, w4_1_18, w4_2_32);
  logic w5_0_7;
  logic w4_2_36;
  csan1 csan4_1_20_4_1_22_X_X_X(w4_1_20, w4_1_22, w4_2_36);
  logic w5_0_8;
  logic w4_2_40;
  csan1 csan4_1_24_4_1_26_X_X_X(w4_1_24, w4_1_26, w4_2_40);
  logic w5_0_9;
  logic w4_3_48;
  csan1 csan4_2_32_4_2_36_X_X_X(w4_2_32, w4_2_36, w4_3_48);
  logic w5_0_10;
  logic w4_4_56;
  csan1 csan4_2_40_4_3_48_X_X_X(w4_2_40, w4_3_48, w4_4_56);
  assign s4 = w4_4_56;
 
 

  assign s = {s4,s3,s2,s1,s0};
end
else if (WIDTH == 32) begin
  assign {w0_0_31, w0_0_30, w0_0_29, w0_0_28, w0_0_27, w0_0_26, w0_0_25, w0_0_24, w0_0_23, w0_0_22, w0_0_21, w0_0_20, w0_0_19, w0_0_18, w0_0_17, w0_0_16, w0_0_15, w0_0_14, w0_0_13, w0_0_12, w0_0_11, w0_0_10, w0_0_9, w0_0_8, w0_0_7, w0_0_6, w0_0_5, w0_0_4, w0_0_3, w0_0_2, w0_0_1, w0_0_0} = a;
  logic w1_0_0;
  logic w0_1_63;
  csan2 csan0_0_31_0_0_30_X_X_X(w0_0_31, w0_0_30, w1_0_0, w0_1_63);
  logic w1_0_1;
  logic w0_1_61;
  csan2 csan0_0_29_0_0_28_X_X_X(w0_0_29, w0_0_28, w1_0_1, w0_1_61);
  logic w1_0_2;
  logic w0_1_59;
  csan2 csan0_0_27_0_0_26_X_X_X(w0_0_27, w0_0_26, w1_0_2, w0_1_59);
  logic w1_0_3;
  logic w0_1_57;
  csan2 csan0_0_25_0_0_24_X_X_X(w0_0_25, w0_0_24, w1_0_3, w0_1_57);
  logic w1_0_4;
  logic w0_1_55;
  csan2 csan0_0_23_0_0_22_X_X_X(w0_0_23, w0_0_22, w1_0_4, w0_1_55);
  logic w1_0_5;
  logic w0_1_53;
  csan2 csan0_0_21_0_0_20_X_X_X(w0_0_21, w0_0_20, w1_0_5, w0_1_53);
  logic w1_0_6;
  logic w0_1_51;
  csan2 csan0_0_19_0_0_18_X_X_X(w0_0_19, w0_0_18, w1_0_6, w0_1_51);
  logic w1_0_7;
  logic w0_1_49;
  csan2 csan0_0_17_0_0_16_X_X_X(w0_0_17, w0_0_16, w1_0_7, w0_1_49);
  logic w1_0_8;
  logic w0_1_47;
  csan2 csan0_0_15_0_0_14_X_X_X(w0_0_15, w0_0_14, w1_0_8, w0_1_47);
  logic w1_0_9;
  logic w0_1_45;
  csan2 csan0_0_13_0_0_12_X_X_X(w0_0_13, w0_0_12, w1_0_9, w0_1_45);
  logic w1_0_10;
  logic w0_1_43;
  csan2 csan0_0_11_0_0_10_X_X_X(w0_0_11, w0_0_10, w1_0_10, w0_1_43);
  logic w1_0_11;
  logic w0_1_41;
  csan2 csan0_0_9_0_0_8_X_X_X(w0_0_9, w0_0_8, w1_0_11, w0_1_41);
  logic w1_0_12;
  logic w0_1_39;
  csan2 csan0_0_7_0_0_6_X_X_X(w0_0_7, w0_0_6, w1_0_12, w0_1_39);
  logic w1_0_13;
  logic w0_1_37;
  csan2 csan0_0_5_0_0_4_X_X_X(w0_0_5, w0_0_4, w1_0_13, w0_1_37);
  logic w1_0_14;
  logic w0_1_35;
  csan2 csan0_0_3_0_0_2_X_X_X(w0_0_3, w0_0_2, w1_0_14, w0_1_35);
  logic w1_0_15;
  logic w0_1_33;
  csan2 csan0_0_1_0_0_0_X_X_X(w0_0_1, w0_0_0, w1_0_15, w0_1_33);
  logic w1_0_16;
  logic w0_2_95;
  csan2 csan0_1_63_0_1_61_X_X_X(w0_1_63, w0_1_61, w1_0_16, w0_2_95);
  logic w1_0_17;
  logic w0_2_91;
  csan2 csan0_1_59_0_1_57_X_X_X(w0_1_59, w0_1_57, w1_0_17, w0_2_91);
  logic w1_0_18;
  logic w0_2_87;
  csan2 csan0_1_55_0_1_53_X_X_X(w0_1_55, w0_1_53, w1_0_18, w0_2_87);
  logic w1_0_19;
  logic w0_2_83;
  csan2 csan0_1_51_0_1_49_X_X_X(w0_1_51, w0_1_49, w1_0_19, w0_2_83);
  logic w1_0_20;
  logic w0_2_79;
  csan2 csan0_1_47_0_1_45_X_X_X(w0_1_47, w0_1_45, w1_0_20, w0_2_79);
  logic w1_0_21;
  logic w0_2_75;
  csan2 csan0_1_43_0_1_41_X_X_X(w0_1_43, w0_1_41, w1_0_21, w0_2_75);
  logic w1_0_22;
  logic w0_2_71;
  csan2 csan0_1_39_0_1_37_X_X_X(w0_1_39, w0_1_37, w1_0_22, w0_2_71);
  logic w1_0_23;
  logic w0_2_67;
  csan2 csan0_1_35_0_1_33_X_X_X(w0_1_35, w0_1_33, w1_0_23, w0_2_67);
  logic w1_0_24;
  logic w0_3_127;
  csan2 csan0_2_95_0_2_91_X_X_X(w0_2_95, w0_2_91, w1_0_24, w0_3_127);
  logic w1_0_25;
  logic w0_3_119;
  csan2 csan0_2_87_0_2_83_X_X_X(w0_2_87, w0_2_83, w1_0_25, w0_3_119);
  logic w1_0_26;
  logic w0_3_111;
  csan2 csan0_2_79_0_2_75_X_X_X(w0_2_79, w0_2_75, w1_0_26, w0_3_111);
  logic w1_0_27;
  logic w0_3_103;
  csan2 csan0_2_71_0_2_67_X_X_X(w0_2_71, w0_2_67, w1_0_27, w0_3_103);
  logic w1_0_28;
  logic w0_4_159;
  csan2 csan0_3_127_0_3_119_X_X_X(w0_3_127, w0_3_119, w1_0_28, w0_4_159);
  logic w1_0_29;
  logic w0_4_143;
  csan2 csan0_3_111_0_3_103_X_X_X(w0_3_111, w0_3_103, w1_0_29, w0_4_143);
  logic w1_0_30;
  logic w0_5_191;
  csan2 csan0_4_159_0_4_143_X_X_X(w0_4_159, w0_4_143, w1_0_30, w0_5_191);
  assign s0 = w0_5_191;
  logic w2_0_0;
  logic w1_1_32;
  csan2 csan1_0_0_1_0_1_X_X_X(w1_0_0, w1_0_1, w2_0_0, w1_1_32);
  logic w2_0_1;
  logic w1_1_34;
  csan2 csan1_0_2_1_0_3_X_X_X(w1_0_2, w1_0_3, w2_0_1, w1_1_34);
  logic w2_0_2;
  logic w1_1_36;
  csan2 csan1_0_4_1_0_5_X_X_X(w1_0_4, w1_0_5, w2_0_2, w1_1_36);
  logic w2_0_3;
  logic w1_1_38;
  csan2 csan1_0_6_1_0_7_X_X_X(w1_0_6, w1_0_7, w2_0_3, w1_1_38);
  logic w2_0_4;
  logic w1_1_40;
  csan2 csan1_0_8_1_0_9_X_X_X(w1_0_8, w1_0_9, w2_0_4, w1_1_40);
  logic w2_0_5;
  logic w1_1_42;
  csan2 csan1_0_10_1_0_11_X_X_X(w1_0_10, w1_0_11, w2_0_5, w1_1_42);
  logic w2_0_6;
  logic w1_1_44;
  csan2 csan1_0_12_1_0_13_X_X_X(w1_0_12, w1_0_13, w2_0_6, w1_1_44);
  logic w2_0_7;
  logic w1_1_46;
  csan2 csan1_0_14_1_0_15_X_X_X(w1_0_14, w1_0_15, w2_0_7, w1_1_46);
  logic w2_0_8;
  logic w1_1_48;
  csan2 csan1_0_16_1_0_17_X_X_X(w1_0_16, w1_0_17, w2_0_8, w1_1_48);
  logic w2_0_9;
  logic w1_1_50;
  csan2 csan1_0_18_1_0_19_X_X_X(w1_0_18, w1_0_19, w2_0_9, w1_1_50);
  logic w2_0_10;
  logic w1_1_52;
  csan2 csan1_0_20_1_0_21_X_X_X(w1_0_20, w1_0_21, w2_0_10, w1_1_52);
  logic w2_0_11;
  logic w1_1_54;
  csan2 csan1_0_22_1_0_23_X_X_X(w1_0_22, w1_0_23, w2_0_11, w1_1_54);
  logic w2_0_12;
  logic w1_1_56;
  csan2 csan1_0_24_1_0_25_X_X_X(w1_0_24, w1_0_25, w2_0_12, w1_1_56);
  logic w2_0_13;
  logic w1_1_58;
  csan2 csan1_0_26_1_0_27_X_X_X(w1_0_26, w1_0_27, w2_0_13, w1_1_58);
  logic w2_0_14;
  logic w1_1_60;
  csan2 csan1_0_28_1_0_29_X_X_X(w1_0_28, w1_0_29, w2_0_14, w1_1_60);
  logic w2_0_15;
  logic w1_2_62;
  csan2 csan1_0_30_1_1_32_X_X_X(w1_0_30, w1_1_32, w2_0_15, w1_2_62);
  logic w2_0_16;
  logic w1_2_66;
  csan2 csan1_1_34_1_1_36_X_X_X(w1_1_34, w1_1_36, w2_0_16, w1_2_66);
  logic w2_0_17;
  logic w1_2_70;
  csan2 csan1_1_38_1_1_40_X_X_X(w1_1_38, w1_1_40, w2_0_17, w1_2_70);
  logic w2_0_18;
  logic w1_2_74;
  csan2 csan1_1_42_1_1_44_X_X_X(w1_1_42, w1_1_44, w2_0_18, w1_2_74);
  logic w2_0_19;
  logic w1_2_78;
  csan2 csan1_1_46_1_1_48_X_X_X(w1_1_46, w1_1_48, w2_0_19, w1_2_78);
  logic w2_0_20;
  logic w1_2_82;
  csan2 csan1_1_50_1_1_52_X_X_X(w1_1_50, w1_1_52, w2_0_20, w1_2_82);
  logic w2_0_21;
  logic w1_2_86;
  csan2 csan1_1_54_1_1_56_X_X_X(w1_1_54, w1_1_56, w2_0_21, w1_2_86);
  logic w2_0_22;
  logic w1_2_90;
  csan2 csan1_1_58_1_1_60_X_X_X(w1_1_58, w1_1_60, w2_0_22, w1_2_90);
  logic w2_0_23;
  logic w1_3_94;
  csan2 csan1_2_62_1_2_66_X_X_X(w1_2_62, w1_2_66, w2_0_23, w1_3_94);
  logic w2_0_24;
  logic w1_3_102;
  csan2 csan1_2_70_1_2_74_X_X_X(w1_2_70, w1_2_74, w2_0_24, w1_3_102);
  logic w2_0_25;
  logic w1_3_110;
  csan2 csan1_2_78_1_2_82_X_X_X(w1_2_78, w1_2_82, w2_0_25, w1_3_110);
  logic w2_0_26;
  logic w1_3_118;
  csan2 csan1_2_86_1_2_90_X_X_X(w1_2_86, w1_2_90, w2_0_26, w1_3_118);
  logic w2_0_27;
  logic w1_4_126;
  csan2 csan1_3_94_1_3_102_X_X_X(w1_3_94, w1_3_102, w2_0_27, w1_4_126);
  logic w2_0_28;
  logic w1_4_142;
  csan2 csan1_3_110_1_3_118_X_X_X(w1_3_110, w1_3_118, w2_0_28, w1_4_142);
  logic w2_0_29;
  logic w1_5_158;
  csan2 csan1_4_126_1_4_142_X_X_X(w1_4_126, w1_4_142, w2_0_29, w1_5_158);
  assign s1 = w1_5_158;
  logic w3_0_0;
  logic w2_1_32;
  csan2 csan2_0_0_2_0_1_X_X_X(w2_0_0, w2_0_1, w3_0_0, w2_1_32);
  logic w3_0_1;
  logic w2_1_34;
  csan2 csan2_0_2_2_0_3_X_X_X(w2_0_2, w2_0_3, w3_0_1, w2_1_34);
  logic w3_0_2;
  logic w2_1_36;
  csan2 csan2_0_4_2_0_5_X_X_X(w2_0_4, w2_0_5, w3_0_2, w2_1_36);
  logic w3_0_3;
  logic w2_1_38;
  csan2 csan2_0_6_2_0_7_X_X_X(w2_0_6, w2_0_7, w3_0_3, w2_1_38);
  logic w3_0_4;
  logic w2_1_40;
  csan2 csan2_0_8_2_0_9_X_X_X(w2_0_8, w2_0_9, w3_0_4, w2_1_40);
  logic w3_0_5;
  logic w2_1_42;
  csan2 csan2_0_10_2_0_11_X_X_X(w2_0_10, w2_0_11, w3_0_5, w2_1_42);
  logic w3_0_6;
  logic w2_1_44;
  csan2 csan2_0_12_2_0_13_X_X_X(w2_0_12, w2_0_13, w3_0_6, w2_1_44);
  logic w3_0_7;
  logic w2_1_46;
  csan2 csan2_0_14_2_0_15_X_X_X(w2_0_14, w2_0_15, w3_0_7, w2_1_46);
  logic w3_0_8;
  logic w2_1_48;
  csan2 csan2_0_16_2_0_17_X_X_X(w2_0_16, w2_0_17, w3_0_8, w2_1_48);
  logic w3_0_9;
  logic w2_1_50;
  csan2 csan2_0_18_2_0_19_X_X_X(w2_0_18, w2_0_19, w3_0_9, w2_1_50);
  logic w3_0_10;
  logic w2_1_52;
  csan2 csan2_0_20_2_0_21_X_X_X(w2_0_20, w2_0_21, w3_0_10, w2_1_52);
  logic w3_0_11;
  logic w2_1_54;
  csan2 csan2_0_22_2_0_23_X_X_X(w2_0_22, w2_0_23, w3_0_11, w2_1_54);
  logic w3_0_12;
  logic w2_1_56;
  csan2 csan2_0_24_2_0_25_X_X_X(w2_0_24, w2_0_25, w3_0_12, w2_1_56);
  logic w3_0_13;
  logic w2_1_58;
  csan2 csan2_0_26_2_0_27_X_X_X(w2_0_26, w2_0_27, w3_0_13, w2_1_58);
  logic w3_0_14;
  logic w2_1_60;
  csan2 csan2_0_28_2_0_29_X_X_X(w2_0_28, w2_0_29, w3_0_14, w2_1_60);
  logic w3_0_15;
  logic w2_2_64;
  csan2 csan2_1_32_2_1_34_X_X_X(w2_1_32, w2_1_34, w3_0_15, w2_2_64);
  logic w3_0_16;
  logic w2_2_68;
  csan2 csan2_1_36_2_1_38_X_X_X(w2_1_36, w2_1_38, w3_0_16, w2_2_68);
  logic w3_0_17;
  logic w2_2_72;
  csan2 csan2_1_40_2_1_42_X_X_X(w2_1_40, w2_1_42, w3_0_17, w2_2_72);
  logic w3_0_18;
  logic w2_2_76;
  csan2 csan2_1_44_2_1_46_X_X_X(w2_1_44, w2_1_46, w3_0_18, w2_2_76);
  logic w3_0_19;
  logic w2_2_80;
  csan2 csan2_1_48_2_1_50_X_X_X(w2_1_48, w2_1_50, w3_0_19, w2_2_80);
  logic w3_0_20;
  logic w2_2_84;
  csan2 csan2_1_52_2_1_54_X_X_X(w2_1_52, w2_1_54, w3_0_20, w2_2_84);
  logic w3_0_21;
  logic w2_2_88;
  csan2 csan2_1_56_2_1_58_X_X_X(w2_1_56, w2_1_58, w3_0_21, w2_2_88);
  logic w3_0_22;
  logic w2_3_92;
  csan2 csan2_1_60_2_2_64_X_X_X(w2_1_60, w2_2_64, w3_0_22, w2_3_92);
  logic w3_0_23;
  logic w2_3_100;
  csan2 csan2_2_68_2_2_72_X_X_X(w2_2_68, w2_2_72, w3_0_23, w2_3_100);
  logic w3_0_24;
  logic w2_3_108;
  csan2 csan2_2_76_2_2_80_X_X_X(w2_2_76, w2_2_80, w3_0_24, w2_3_108);
  logic w3_0_25;
  logic w2_3_116;
  csan2 csan2_2_84_2_2_88_X_X_X(w2_2_84, w2_2_88, w3_0_25, w2_3_116);
  logic w3_0_26;
  logic w2_4_124;
  csan2 csan2_3_92_2_3_100_X_X_X(w2_3_92, w2_3_100, w3_0_26, w2_4_124);
  logic w3_0_27;
  logic w2_4_140;
  csan2 csan2_3_108_2_3_116_X_X_X(w2_3_108, w2_3_116, w3_0_27, w2_4_140);
  logic w3_0_28;
  logic w2_5_156;
  csan2 csan2_4_124_2_4_140_X_X_X(w2_4_124, w2_4_140, w3_0_28, w2_5_156);
  assign s2 = w2_5_156;
  logic w4_0_0;
  logic w3_1_32;
  csan2 csan3_0_0_3_0_1_X_X_X(w3_0_0, w3_0_1, w4_0_0, w3_1_32);
  logic w4_0_1;
  logic w3_1_34;
  csan2 csan3_0_2_3_0_3_X_X_X(w3_0_2, w3_0_3, w4_0_1, w3_1_34);
  logic w4_0_2;
  logic w3_1_36;
  csan2 csan3_0_4_3_0_5_X_X_X(w3_0_4, w3_0_5, w4_0_2, w3_1_36);
  logic w4_0_3;
  logic w3_1_38;
  csan2 csan3_0_6_3_0_7_X_X_X(w3_0_6, w3_0_7, w4_0_3, w3_1_38);
  logic w4_0_4;
  logic w3_1_40;
  csan2 csan3_0_8_3_0_9_X_X_X(w3_0_8, w3_0_9, w4_0_4, w3_1_40);
  logic w4_0_5;
  logic w3_1_42;
  csan2 csan3_0_10_3_0_11_X_X_X(w3_0_10, w3_0_11, w4_0_5, w3_1_42);
  logic w4_0_6;
  logic w3_1_44;
  csan2 csan3_0_12_3_0_13_X_X_X(w3_0_12, w3_0_13, w4_0_6, w3_1_44);
  logic w4_0_7;
  logic w3_1_46;
  csan2 csan3_0_14_3_0_15_X_X_X(w3_0_14, w3_0_15, w4_0_7, w3_1_46);
  logic w4_0_8;
  logic w3_1_48;
  csan2 csan3_0_16_3_0_17_X_X_X(w3_0_16, w3_0_17, w4_0_8, w3_1_48);
  logic w4_0_9;
  logic w3_1_50;
  csan2 csan3_0_18_3_0_19_X_X_X(w3_0_18, w3_0_19, w4_0_9, w3_1_50);
  logic w4_0_10;
  logic w3_1_52;
  csan2 csan3_0_20_3_0_21_X_X_X(w3_0_20, w3_0_21, w4_0_10, w3_1_52);
  logic w4_0_11;
  logic w3_1_54;
  csan2 csan3_0_22_3_0_23_X_X_X(w3_0_22, w3_0_23, w4_0_11, w3_1_54);
  logic w4_0_12;
  logic w3_1_56;
  csan2 csan3_0_24_3_0_25_X_X_X(w3_0_24, w3_0_25, w4_0_12, w3_1_56);
  logic w4_0_13;
  logic w3_1_58;
  csan2 csan3_0_26_3_0_27_X_X_X(w3_0_26, w3_0_27, w4_0_13, w3_1_58);
  logic w4_0_14;
  logic w3_2_60;
  csan2 csan3_0_28_3_1_32_X_X_X(w3_0_28, w3_1_32, w4_0_14, w3_2_60);
  logic w4_0_15;
  logic w3_2_66;
  csan2 csan3_1_34_3_1_36_X_X_X(w3_1_34, w3_1_36, w4_0_15, w3_2_66);
  logic w4_0_16;
  logic w3_2_70;
  csan2 csan3_1_38_3_1_40_X_X_X(w3_1_38, w3_1_40, w4_0_16, w3_2_70);
  logic w4_0_17;
  logic w3_2_74;
  csan2 csan3_1_42_3_1_44_X_X_X(w3_1_42, w3_1_44, w4_0_17, w3_2_74);
  logic w4_0_18;
  logic w3_2_78;
  csan2 csan3_1_46_3_1_48_X_X_X(w3_1_46, w3_1_48, w4_0_18, w3_2_78);
  logic w4_0_19;
  logic w3_2_82;
  csan2 csan3_1_50_3_1_52_X_X_X(w3_1_50, w3_1_52, w4_0_19, w3_2_82);
  logic w4_0_20;
  logic w3_2_86;
  csan2 csan3_1_54_3_1_56_X_X_X(w3_1_54, w3_1_56, w4_0_20, w3_2_86);
  logic w4_0_21;
  logic w3_3_90;
  csan2 csan3_1_58_3_2_60_X_X_X(w3_1_58, w3_2_60, w4_0_21, w3_3_90);
  logic w4_0_22;
  logic w3_3_98;
  csan2 csan3_2_66_3_2_70_X_X_X(w3_2_66, w3_2_70, w4_0_22, w3_3_98);
  logic w4_0_23;
  logic w3_3_106;
  csan2 csan3_2_74_3_2_78_X_X_X(w3_2_74, w3_2_78, w4_0_23, w3_3_106);
  logic w4_0_24;
  logic w3_3_114;
  csan2 csan3_2_82_3_2_86_X_X_X(w3_2_82, w3_2_86, w4_0_24, w3_3_114);
  logic w4_0_25;
  logic w3_4_122;
  csan2 csan3_3_90_3_3_98_X_X_X(w3_3_90, w3_3_98, w4_0_25, w3_4_122);
  logic w4_0_26;
  logic w3_4_138;
  csan2 csan3_3_106_3_3_114_X_X_X(w3_3_106, w3_3_114, w4_0_26, w3_4_138);
  logic w4_0_27;
  logic w3_5_154;
  csan2 csan3_4_122_3_4_138_X_X_X(w3_4_122, w3_4_138, w4_0_27, w3_5_154);
  assign s3 = w3_5_154;
  logic w5_0_0;
  logic w4_1_32;
  csan2 csan4_0_0_4_0_1_X_X_X(w4_0_0, w4_0_1, w5_0_0, w4_1_32);
  logic w5_0_1;
  logic w4_1_34;
  csan2 csan4_0_2_4_0_3_X_X_X(w4_0_2, w4_0_3, w5_0_1, w4_1_34);
  logic w5_0_2;
  logic w4_1_36;
  csan2 csan4_0_4_4_0_5_X_X_X(w4_0_4, w4_0_5, w5_0_2, w4_1_36);
  logic w5_0_3;
  logic w4_1_38;
  csan2 csan4_0_6_4_0_7_X_X_X(w4_0_6, w4_0_7, w5_0_3, w4_1_38);
  logic w5_0_4;
  logic w4_1_40;
  csan2 csan4_0_8_4_0_9_X_X_X(w4_0_8, w4_0_9, w5_0_4, w4_1_40);
  logic w5_0_5;
  logic w4_1_42;
  csan2 csan4_0_10_4_0_11_X_X_X(w4_0_10, w4_0_11, w5_0_5, w4_1_42);
  logic w5_0_6;
  logic w4_1_44;
  csan2 csan4_0_12_4_0_13_X_X_X(w4_0_12, w4_0_13, w5_0_6, w4_1_44);
  logic w5_0_7;
  logic w4_1_46;
  csan2 csan4_0_14_4_0_15_X_X_X(w4_0_14, w4_0_15, w5_0_7, w4_1_46);
  logic w5_0_8;
  logic w4_1_48;
  csan2 csan4_0_16_4_0_17_X_X_X(w4_0_16, w4_0_17, w5_0_8, w4_1_48);
  logic w5_0_9;
  logic w4_1_50;
  csan2 csan4_0_18_4_0_19_X_X_X(w4_0_18, w4_0_19, w5_0_9, w4_1_50);
  logic w5_0_10;
  logic w4_1_52;
  csan2 csan4_0_20_4_0_21_X_X_X(w4_0_20, w4_0_21, w5_0_10, w4_1_52);
  logic w5_0_11;
  logic w4_1_54;
  csan2 csan4_0_22_4_0_23_X_X_X(w4_0_22, w4_0_23, w5_0_11, w4_1_54);
  logic w5_0_12;
  logic w4_1_56;
  csan2 csan4_0_24_4_0_25_X_X_X(w4_0_24, w4_0_25, w5_0_12, w4_1_56);
  logic w5_0_13;
  logic w4_1_58;
  csan2 csan4_0_26_4_0_27_X_X_X(w4_0_26, w4_0_27, w5_0_13, w4_1_58);
  logic w5_0_14;
  logic w4_2_64;
  csan2 csan4_1_32_4_1_34_X_X_X(w4_1_32, w4_1_34, w5_0_14, w4_2_64);
  logic w5_0_15;
  logic w4_2_68;
  csan2 csan4_1_36_4_1_38_X_X_X(w4_1_36, w4_1_38, w5_0_15, w4_2_68);
  logic w5_0_16;
  logic w4_2_72;
  csan2 csan4_1_40_4_1_42_X_X_X(w4_1_40, w4_1_42, w5_0_16, w4_2_72);
  logic w5_0_17;
  logic w4_2_76;
  csan2 csan4_1_44_4_1_46_X_X_X(w4_1_44, w4_1_46, w5_0_17, w4_2_76);
  logic w5_0_18;
  logic w4_2_80;
  csan2 csan4_1_48_4_1_50_X_X_X(w4_1_48, w4_1_50, w5_0_18, w4_2_80);
  logic w5_0_19;
  logic w4_2_84;
  csan2 csan4_1_52_4_1_54_X_X_X(w4_1_52, w4_1_54, w5_0_19, w4_2_84);
  logic w5_0_20;
  logic w4_2_88;
  csan2 csan4_1_56_4_1_58_X_X_X(w4_1_56, w4_1_58, w5_0_20, w4_2_88);
  logic w5_0_21;
  logic w4_3_96;
  csan2 csan4_2_64_4_2_68_X_X_X(w4_2_64, w4_2_68, w5_0_21, w4_3_96);
  logic w5_0_22;
  logic w4_3_104;
  csan2 csan4_2_72_4_2_76_X_X_X(w4_2_72, w4_2_76, w5_0_22, w4_3_104);
  logic w5_0_23;
  logic w4_3_112;
  csan2 csan4_2_80_4_2_84_X_X_X(w4_2_80, w4_2_84, w5_0_23, w4_3_112);
  logic w5_0_24;
  logic w4_4_120;
  csan2 csan4_2_88_4_3_96_X_X_X(w4_2_88, w4_3_96, w5_0_24, w4_4_120);
  logic w5_0_25;
  logic w4_4_136;
  csan2 csan4_3_104_4_3_112_X_X_X(w4_3_104, w4_3_112, w5_0_25, w4_4_136);
  logic w5_0_26;
  logic w4_5_152;
  csan2 csan4_4_120_4_4_136_X_X_X(w4_4_120, w4_4_136, w5_0_26, w4_5_152);
  assign s4 = w4_5_152;
  logic w6_0_0;
  logic w5_1_32;
  csan2 csan5_0_0_5_0_1_X_X_X(w5_0_0, w5_0_1, w6_0_0, w5_1_32);
  logic w6_0_1;
  logic w5_1_34;
  csan2 csan5_0_2_5_0_3_X_X_X(w5_0_2, w5_0_3, w6_0_1, w5_1_34);
  logic w6_0_2;
  logic w5_1_36;
  csan2 csan5_0_4_5_0_5_X_X_X(w5_0_4, w5_0_5, w6_0_2, w5_1_36);
  logic w6_0_3;
  logic w5_1_38;
  csan2 csan5_0_6_5_0_7_X_X_X(w5_0_6, w5_0_7, w6_0_3, w5_1_38);
  logic w6_0_4;
  logic w5_1_40;
  csan2 csan5_0_8_5_0_9_X_X_X(w5_0_8, w5_0_9, w6_0_4, w5_1_40);
  logic w6_0_5;
  logic w5_1_42;
  csan2 csan5_0_10_5_0_11_X_X_X(w5_0_10, w5_0_11, w6_0_5, w5_1_42);
  logic w6_0_6;
  logic w5_1_44;
  csan2 csan5_0_12_5_0_13_X_X_X(w5_0_12, w5_0_13, w6_0_6, w5_1_44);
  logic w6_0_7;
  logic w5_1_46;
  csan2 csan5_0_14_5_0_15_X_X_X(w5_0_14, w5_0_15, w6_0_7, w5_1_46);
  logic w6_0_8;
  logic w5_1_48;
  csan2 csan5_0_16_5_0_17_X_X_X(w5_0_16, w5_0_17, w6_0_8, w5_1_48);
  logic w6_0_9;
  logic w5_1_50;
  csan2 csan5_0_18_5_0_19_X_X_X(w5_0_18, w5_0_19, w6_0_9, w5_1_50);
  logic w6_0_10;
  logic w5_1_52;
  csan2 csan5_0_20_5_0_21_X_X_X(w5_0_20, w5_0_21, w6_0_10, w5_1_52);
  logic w6_0_11;
  logic w5_1_54;
  csan2 csan5_0_22_5_0_23_X_X_X(w5_0_22, w5_0_23, w6_0_11, w5_1_54);
  logic w6_0_12;
  logic w5_1_56;
  csan2 csan5_0_24_5_0_25_X_X_X(w5_0_24, w5_0_25, w6_0_12, w5_1_56);
  logic w6_0_13;
  logic w5_2_58;
  csan2 csan5_0_26_5_1_32_X_X_X(w5_0_26, w5_1_32, w6_0_13, w5_2_58);
  logic w6_0_14;
  logic w5_2_66;
  csan2 csan5_1_34_5_1_36_X_X_X(w5_1_34, w5_1_36, w6_0_14, w5_2_66);
  logic w6_0_15;
  logic w5_2_70;
  csan2 csan5_1_38_5_1_40_X_X_X(w5_1_38, w5_1_40, w6_0_15, w5_2_70);
  logic w6_0_16;
  logic w5_2_74;
  csan2 csan5_1_42_5_1_44_X_X_X(w5_1_42, w5_1_44, w6_0_16, w5_2_74);
  logic w6_0_17;
  logic w5_2_78;
  csan2 csan5_1_46_5_1_48_X_X_X(w5_1_46, w5_1_48, w6_0_17, w5_2_78);
  logic w6_0_18;
  logic w5_2_82;
  csan2 csan5_1_50_5_1_52_X_X_X(w5_1_50, w5_1_52, w6_0_18, w5_2_82);
  logic w6_0_19;
  logic w5_2_86;
  csan2 csan5_1_54_5_1_56_X_X_X(w5_1_54, w5_1_56, w6_0_19, w5_2_86);
  logic w6_0_20;
  logic w5_3_90;
  csan2 csan5_2_58_5_2_66_X_X_X(w5_2_58, w5_2_66, w6_0_20, w5_3_90);
  logic w6_0_21;
  logic w5_3_102;
  csan2 csan5_2_70_5_2_74_X_X_X(w5_2_70, w5_2_74, w6_0_21, w5_3_102);
  logic w6_0_22;
  logic w5_3_110;
  csan2 csan5_2_78_5_2_82_X_X_X(w5_2_78, w5_2_82, w6_0_22, w5_3_110);
  logic w6_0_23;
  logic w5_4_118;
  csan2 csan5_2_86_5_3_90_X_X_X(w5_2_86, w5_3_90, w6_0_23, w5_4_118);
  logic w6_0_24;
  logic w5_4_134;
  csan2 csan5_3_102_5_3_110_X_X_X(w5_3_102, w5_3_110, w6_0_24, w5_4_134);
  logic w6_0_25;
  logic w5_5_150;
  csan2 csan5_4_118_5_4_134_X_X_X(w5_4_118, w5_4_134, w6_0_25, w5_5_150);
  assign s5 = w5_5_150;
  assign s = {s5, s4, s3, s2, s1, s0};
end else begin

  assign {w0_0_63, w0_0_62, w0_0_61, w0_0_60, w0_0_59, w0_0_58, w0_0_57, w0_0_56, w0_0_55, w0_0_54, w0_0_53, w0_0_52, w0_0_51, w0_0_50, w0_0_49, w0_0_48, w0_0_47, w0_0_46, w0_0_45, w0_0_44, w0_0_43, w0_0_42, w0_0_41, w0_0_40, w0_0_39, w0_0_38, w0_0_37, w0_0_36, w0_0_35, w0_0_34, w0_0_33, w0_0_32, w0_0_31, w0_0_30, w0_0_29, w0_0_28, w0_0_27, w0_0_26, w0_0_25, w0_0_24, w0_0_23, w0_0_22, w0_0_21, w0_0_20, w0_0_19, w0_0_18, w0_0_17, w0_0_16, w0_0_15, w0_0_14, w0_0_13, w0_0_12, w0_0_11, w0_0_10, w0_0_9, w0_0_8, w0_0_7, w0_0_6, w0_0_5, w0_0_4, w0_0_3, w0_0_2, w0_0_1, w0_0_0} = a;
  logic w1_0_0;
  logic w0_1_127;
  csan csan0_0_63_0_0_62_0_0_61(w0_0_63, w0_0_62, w0_0_61, w1_0_0, w0_1_127);
  logic w1_0_1;
  logic w0_1_124;
  csan csan0_0_60_0_0_59_0_0_58(w0_0_60, w0_0_59, w0_0_58, w1_0_1, w0_1_124);
  logic w1_0_2;
  logic w0_1_121;
  csan csan0_0_57_0_0_56_0_0_55(w0_0_57, w0_0_56, w0_0_55, w1_0_2, w0_1_121);
  logic w1_0_3;
  logic w0_1_118;
  csan csan0_0_54_0_0_53_0_0_52(w0_0_54, w0_0_53, w0_0_52, w1_0_3, w0_1_118);
  logic w1_0_4;
  logic w0_1_115;
  csan csan0_0_51_0_0_50_0_0_49(w0_0_51, w0_0_50, w0_0_49, w1_0_4, w0_1_115);
  logic w1_0_5;
  logic w0_1_112;
  csan csan0_0_48_0_0_47_0_0_46(w0_0_48, w0_0_47, w0_0_46, w1_0_5, w0_1_112);
  logic w1_0_6;
  logic w0_1_109;
  csan csan0_0_45_0_0_44_0_0_43(w0_0_45, w0_0_44, w0_0_43, w1_0_6, w0_1_109);
  logic w1_0_7;
  logic w0_1_106;
  csan csan0_0_42_0_0_41_0_0_40(w0_0_42, w0_0_41, w0_0_40, w1_0_7, w0_1_106);
  logic w1_0_8;
  logic w0_1_103;
  csan csan0_0_39_0_0_38_0_0_37(w0_0_39, w0_0_38, w0_0_37, w1_0_8, w0_1_103);
  logic w1_0_9;
  logic w0_1_100;
  csan csan0_0_36_0_0_35_0_0_34(w0_0_36, w0_0_35, w0_0_34, w1_0_9, w0_1_100);
  logic w1_0_10;
  logic w0_1_97;
  csan csan0_0_33_0_0_32_0_0_31(w0_0_33, w0_0_32, w0_0_31, w1_0_10, w0_1_97);
  logic w1_0_11;
  logic w0_1_94;
  csan csan0_0_30_0_0_29_0_0_28(w0_0_30, w0_0_29, w0_0_28, w1_0_11, w0_1_94);
  logic w1_0_12;
  logic w0_1_91;
  csan csan0_0_27_0_0_26_0_0_25(w0_0_27, w0_0_26, w0_0_25, w1_0_12, w0_1_91);
  logic w1_0_13;
  logic w0_1_88;
  csan csan0_0_24_0_0_23_0_0_22(w0_0_24, w0_0_23, w0_0_22, w1_0_13, w0_1_88);
  logic w1_0_14;
  logic w0_1_85;
  csan csan0_0_21_0_0_20_0_0_19(w0_0_21, w0_0_20, w0_0_19, w1_0_14, w0_1_85);
  logic w1_0_15;
  logic w0_1_82;
  csan csan0_0_18_0_0_17_0_0_16(w0_0_18, w0_0_17, w0_0_16, w1_0_15, w0_1_82);
  logic w1_0_16;
  logic w0_1_79;
  csan csan0_0_15_0_0_14_0_0_13(w0_0_15, w0_0_14, w0_0_13, w1_0_16, w0_1_79);
  logic w1_0_17;
  logic w0_1_76;
  csan csan0_0_12_0_0_11_0_0_10(w0_0_12, w0_0_11, w0_0_10, w1_0_17, w0_1_76);
  logic w1_0_18;
  logic w0_1_73;
  csan csan0_0_9_0_0_8_0_0_7(w0_0_9, w0_0_8, w0_0_7, w1_0_18, w0_1_73);
  logic w1_0_19;
  logic w0_1_70;
  csan csan0_0_6_0_0_5_0_0_4(w0_0_6, w0_0_5, w0_0_4, w1_0_19, w0_1_70);
  logic w1_0_20;
  logic w0_1_67;
  csan csan0_0_3_0_0_2_0_0_1(w0_0_3, w0_0_2, w0_0_1, w1_0_20, w0_1_67);
  logic w1_0_21;
  logic w0_2_64;
  csan csan0_0_0_0_1_127_0_1_124(w0_0_0, w0_1_127, w0_1_124, w1_0_21, w0_2_64);
  logic w1_0_22;
  logic w0_2_185;
  csan csan0_1_121_0_1_118_0_1_115(w0_1_121, w0_1_118, w0_1_115, w1_0_22, w0_2_185);
  logic w1_0_23;
  logic w0_2_176;
  csan csan0_1_112_0_1_109_0_1_106(w0_1_112, w0_1_109, w0_1_106, w1_0_23, w0_2_176);
  logic w1_0_24;
  logic w0_2_167;
  csan csan0_1_103_0_1_100_0_1_97(w0_1_103, w0_1_100, w0_1_97, w1_0_24, w0_2_167);
  logic w1_0_25;
  logic w0_2_158;
  csan csan0_1_94_0_1_91_0_1_88(w0_1_94, w0_1_91, w0_1_88, w1_0_25, w0_2_158);
  logic w1_0_26;
  logic w0_2_149;
  csan csan0_1_85_0_1_82_0_1_79(w0_1_85, w0_1_82, w0_1_79, w1_0_26, w0_2_149);
  logic w1_0_27;
  logic w0_2_140;
  csan csan0_1_76_0_1_73_0_1_70(w0_1_76, w0_1_73, w0_1_70, w1_0_27, w0_2_140);
  logic w1_0_28;
  logic w0_3_131;
  csan csan0_1_67_0_2_64_0_2_185(w0_1_67, w0_2_64, w0_2_185, w1_0_28, w0_3_131);
  logic w1_0_29;
  logic w0_3_240;
  csan csan0_2_176_0_2_167_0_2_158(w0_2_176, w0_2_167, w0_2_158, w1_0_29, w0_3_240);
  logic w1_0_30;
  logic w0_4_213;
  csan csan0_2_149_0_2_140_0_3_131(w0_2_149, w0_2_140, w0_3_131, w1_0_30, w0_4_213);
  logic w1_0_31;
  logic w0_5_304;
  csan2 csan0_3_240_0_4_213_X_X_X(w0_3_240, w0_4_213, w1_0_31, w0_5_304);
  assign s0 = w0_5_304;
  logic w2_0_0;
  logic w1_1_64;
  csan csan1_0_0_1_0_1_1_0_2(w1_0_0, w1_0_1, w1_0_2, w2_0_0, w1_1_64);
  logic w2_0_1;
  logic w1_1_67;
  csan csan1_0_3_1_0_4_1_0_5(w1_0_3, w1_0_4, w1_0_5, w2_0_1, w1_1_67);
  logic w2_0_2;
  logic w1_1_70;
  csan csan1_0_6_1_0_7_1_0_8(w1_0_6, w1_0_7, w1_0_8, w2_0_2, w1_1_70);
  logic w2_0_3;
  logic w1_1_73;
  csan csan1_0_9_1_0_10_1_0_11(w1_0_9, w1_0_10, w1_0_11, w2_0_3, w1_1_73);
  logic w2_0_4;
  logic w1_1_76;
  csan csan1_0_12_1_0_13_1_0_14(w1_0_12, w1_0_13, w1_0_14, w2_0_4, w1_1_76);
  logic w2_0_5;
  logic w1_1_79;
  csan csan1_0_15_1_0_16_1_0_17(w1_0_15, w1_0_16, w1_0_17, w2_0_5, w1_1_79);
  logic w2_0_6;
  logic w1_1_82;
  csan csan1_0_18_1_0_19_1_0_20(w1_0_18, w1_0_19, w1_0_20, w2_0_6, w1_1_82);
  logic w2_0_7;
  logic w1_1_85;
  csan csan1_0_21_1_0_22_1_0_23(w1_0_21, w1_0_22, w1_0_23, w2_0_7, w1_1_85);
  logic w2_0_8;
  logic w1_1_88;
  csan csan1_0_24_1_0_25_1_0_26(w1_0_24, w1_0_25, w1_0_26, w2_0_8, w1_1_88);
  logic w2_0_9;
  logic w1_1_91;
  csan csan1_0_27_1_0_28_1_0_29(w1_0_27, w1_0_28, w1_0_29, w2_0_9, w1_1_91);
  logic w2_0_10;
  logic w1_2_94;
  csan csan1_0_30_1_0_31_1_1_64(w1_0_30, w1_0_31, w1_1_64, w2_0_10, w1_2_94);
  logic w2_0_11;
  logic w1_2_131;
  csan csan1_1_67_1_1_70_1_1_73(w1_1_67, w1_1_70, w1_1_73, w2_0_11, w1_2_131);
  logic w2_0_12;
  logic w1_2_140;
  csan csan1_1_76_1_1_79_1_1_82(w1_1_76, w1_1_79, w1_1_82, w2_0_12, w1_2_140);
  logic w2_0_13;
  logic w1_2_149;
  csan csan1_1_85_1_1_88_1_1_91(w1_1_85, w1_1_88, w1_1_91, w2_0_13, w1_2_149);
  logic w2_0_14;
  logic w1_3_158;
  csan csan1_2_94_1_2_131_1_2_140(w1_2_94, w1_2_131, w1_2_140, w2_0_14, w1_3_158);
  logic w2_0_15;
  logic w1_4_213;
  csan2 csan1_2_149_1_3_158_X_X_X(w1_2_149, w1_3_158, w2_0_15, w1_4_213);
  assign s1 = w1_4_213;
  logic w3_0_0;
  logic w2_1_64;
  csan csan2_0_0_2_0_1_2_0_2(w2_0_0, w2_0_1, w2_0_2, w3_0_0, w2_1_64);
  logic w3_0_1;
  logic w2_1_67;
  csan csan2_0_3_2_0_4_2_0_5(w2_0_3, w2_0_4, w2_0_5, w3_0_1, w2_1_67);
  logic w3_0_2;
  logic w2_1_70;
  csan csan2_0_6_2_0_7_2_0_8(w2_0_6, w2_0_7, w2_0_8, w3_0_2, w2_1_70);
  logic w3_0_3;
  logic w2_1_73;
  csan csan2_0_9_2_0_10_2_0_11(w2_0_9, w2_0_10, w2_0_11, w3_0_3, w2_1_73);
  logic w3_0_4;
  logic w2_1_76;
  csan csan2_0_12_2_0_13_2_0_14(w2_0_12, w2_0_13, w2_0_14, w3_0_4, w2_1_76);
  logic w3_0_5;
  logic w2_2_79;
  csan csan2_0_15_2_1_64_2_1_67(w2_0_15, w2_1_64, w2_1_67, w3_0_5, w2_2_79);
  logic w3_0_6;
  logic w2_2_134;
  csan csan2_1_70_2_1_73_2_1_76(w2_1_70, w2_1_73, w2_1_76, w3_0_6, w2_2_134);
  logic w3_0_7;
  logic w2_3_143;
  csan2 csan2_2_79_2_2_134_X_X_X(w2_2_79, w2_2_134, w3_0_7, w2_3_143);
  assign s2 = w2_3_143;
  logic w4_0_0;
  logic w3_1_64;
  csan csan3_0_0_3_0_1_3_0_2(w3_0_0, w3_0_1, w3_0_2, w4_0_0, w3_1_64);
  logic w4_0_1;
  logic w3_1_67;
  csan csan3_0_3_3_0_4_3_0_5(w3_0_3, w3_0_4, w3_0_5, w4_0_1, w3_1_67);
  logic w4_0_2;
  logic w3_2_70;
  csan csan3_0_6_3_0_7_3_1_64(w3_0_6, w3_0_7, w3_1_64, w4_0_2, w3_2_70);
  logic w4_0_3;
  logic w3_3_131;
  csan2 csan3_1_67_3_2_70_X_X_X(w3_1_67, w3_2_70, w4_0_3, w3_3_131);
  assign s3 = w3_3_131;
  logic w5_0_0;
  logic w4_1_64;
  csan csan4_0_0_4_0_1_4_0_2(w4_0_0, w4_0_1, w4_0_2, w5_0_0, w4_1_64);
  logic w5_0_1;
  logic w4_2_67;
  csan2 csan4_0_3_4_1_64_X_X_X(w4_0_3, w4_1_64, w5_0_1, w4_2_67);
  assign s4 = w4_2_67;
  logic w6_0_0;
  logic w5_1_64;
  csan2 csan5_0_0_5_0_1_X_X_X(w5_0_0, w5_0_1, w6_0_0, w5_1_64);
  assign s5 = w5_1_64;
  assign s6 = w6_0_0;
  assign s = {s6,s5, s4, s3, s2, s1, s0};
end

endmodule